module Reorder_Buffer(
  input         clock,
  input         reset,
  output        io_o_full,
  input         io_i_rob_allocation_reqs_0_valid,
  input  [31:0] io_i_rob_allocation_reqs_0_uop_pc,
  input  [31:0] io_i_rob_allocation_reqs_0_uop_inst,
  input  [6:0]  io_i_rob_allocation_reqs_0_uop_func_code,
  input  [6:0]  io_i_rob_allocation_reqs_0_uop_phy_dst,
  input  [6:0]  io_i_rob_allocation_reqs_0_uop_stale_dst,
  input  [4:0]  io_i_rob_allocation_reqs_0_uop_arch_dst,
  input  [63:0] io_i_rob_allocation_reqs_0_uop_src1_value,
  input  [4:0]  io_i_rob_allocation_reqs_0_uop_alu_sel,
  input         io_i_rob_allocation_reqs_1_valid,
  input  [31:0] io_i_rob_allocation_reqs_1_uop_pc,
  input  [31:0] io_i_rob_allocation_reqs_1_uop_inst,
  input  [6:0]  io_i_rob_allocation_reqs_1_uop_func_code,
  input  [6:0]  io_i_rob_allocation_reqs_1_uop_phy_dst,
  input  [6:0]  io_i_rob_allocation_reqs_1_uop_stale_dst,
  input  [4:0]  io_i_rob_allocation_reqs_1_uop_arch_dst,
  input  [63:0] io_i_rob_allocation_reqs_1_uop_src1_value,
  input  [4:0]  io_i_rob_allocation_reqs_1_uop_alu_sel,
  output [6:0]  io_o_rob_allocation_ress_0_rob_idx,
  output [6:0]  io_o_rob_allocation_ress_1_rob_idx,
  output        io_o_rollback_packs_0_valid,
  output [6:0]  io_o_rollback_packs_0_uop_phy_dst,
  output [6:0]  io_o_rollback_packs_0_uop_stale_dst,
  output [4:0]  io_o_rollback_packs_0_uop_arch_dst,
  output        io_o_rollback_packs_1_valid,
  output [6:0]  io_o_rollback_packs_1_uop_phy_dst,
  output [6:0]  io_o_rollback_packs_1_uop_stale_dst,
  output [4:0]  io_o_rollback_packs_1_uop_arch_dst,
  input         io_i_ex_res_packs_0_valid,
  input  [31:0] io_i_ex_res_packs_0_uop_pc,
  input  [31:0] io_i_ex_res_packs_0_uop_inst,
  input  [6:0]  io_i_ex_res_packs_0_uop_func_code,
  input  [6:0]  io_i_ex_res_packs_0_uop_phy_dst,
  input  [6:0]  io_i_ex_res_packs_0_uop_stale_dst,
  input  [4:0]  io_i_ex_res_packs_0_uop_arch_dst,
  input  [6:0]  io_i_ex_res_packs_0_uop_rob_idx,
  input  [63:0] io_i_ex_res_packs_0_uop_dst_value,
  input  [63:0] io_i_ex_res_packs_0_uop_src1_value,
  input  [4:0]  io_i_ex_res_packs_0_uop_alu_sel,
  input         io_i_ex_res_packs_1_valid,
  input  [31:0] io_i_ex_res_packs_1_uop_pc,
  input  [31:0] io_i_ex_res_packs_1_uop_inst,
  input  [6:0]  io_i_ex_res_packs_1_uop_func_code,
  input  [6:0]  io_i_ex_res_packs_1_uop_phy_dst,
  input  [6:0]  io_i_ex_res_packs_1_uop_stale_dst,
  input  [4:0]  io_i_ex_res_packs_1_uop_arch_dst,
  input  [6:0]  io_i_ex_res_packs_1_uop_rob_idx,
  input  [63:0] io_i_ex_res_packs_1_uop_dst_value,
  input  [63:0] io_i_ex_res_packs_1_uop_src1_value,
  input  [4:0]  io_i_ex_res_packs_1_uop_alu_sel,
  input         io_i_branch_resolve_pack_valid,
  input         io_i_branch_resolve_pack_mispred,
  input  [7:0]  io_i_branch_resolve_pack_rob_idx,
  output        io_o_commit_packs_0_valid,
  output [31:0] io_o_commit_packs_0_uop_pc,
  output [31:0] io_o_commit_packs_0_uop_inst,
  output [6:0]  io_o_commit_packs_0_uop_func_code,
  output [6:0]  io_o_commit_packs_0_uop_phy_dst,
  output [6:0]  io_o_commit_packs_0_uop_stale_dst,
  output [4:0]  io_o_commit_packs_0_uop_arch_dst,
  output [63:0] io_o_commit_packs_0_uop_dst_value,
  output [63:0] io_o_commit_packs_0_uop_src1_value,
  output [4:0]  io_o_commit_packs_0_uop_alu_sel,
  output        io_o_commit_packs_1_valid,
  output [31:0] io_o_commit_packs_1_uop_inst,
  output [6:0]  io_o_commit_packs_1_uop_func_code,
  output [6:0]  io_o_commit_packs_1_uop_phy_dst,
  output [6:0]  io_o_commit_packs_1_uop_stale_dst,
  output [4:0]  io_o_commit_packs_1_uop_arch_dst,
  output [63:0] io_o_commit_packs_1_uop_dst_value,
  output [63:0] io_o_commit_packs_1_uop_src1_value,
  output [4:0]  io_o_commit_packs_1_uop_alu_sel,
  output [6:0]  io_o_rob_head,
  input         io_i_interrupt,
  input         io_i_csr_pc_redirect,
  output        io_o_exception
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [63:0] _RAND_75;
  reg [63:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [63:0] _RAND_84;
  reg [63:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [63:0] _RAND_93;
  reg [63:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [63:0] _RAND_102;
  reg [63:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [63:0] _RAND_111;
  reg [63:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [63:0] _RAND_120;
  reg [63:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [63:0] _RAND_129;
  reg [63:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [63:0] _RAND_138;
  reg [63:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [63:0] _RAND_147;
  reg [63:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [63:0] _RAND_156;
  reg [63:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [63:0] _RAND_165;
  reg [63:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [63:0] _RAND_174;
  reg [63:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [63:0] _RAND_183;
  reg [63:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [63:0] _RAND_192;
  reg [63:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [63:0] _RAND_201;
  reg [63:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [63:0] _RAND_210;
  reg [63:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [63:0] _RAND_219;
  reg [63:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [63:0] _RAND_228;
  reg [63:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [63:0] _RAND_237;
  reg [63:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [63:0] _RAND_246;
  reg [63:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [63:0] _RAND_255;
  reg [63:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [63:0] _RAND_264;
  reg [63:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [63:0] _RAND_273;
  reg [63:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [63:0] _RAND_282;
  reg [63:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [63:0] _RAND_291;
  reg [63:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [63:0] _RAND_300;
  reg [63:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [63:0] _RAND_309;
  reg [63:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [63:0] _RAND_318;
  reg [63:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [63:0] _RAND_327;
  reg [63:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [63:0] _RAND_336;
  reg [63:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [63:0] _RAND_345;
  reg [63:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [63:0] _RAND_354;
  reg [63:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [63:0] _RAND_363;
  reg [63:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [63:0] _RAND_372;
  reg [63:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [63:0] _RAND_381;
  reg [63:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [63:0] _RAND_390;
  reg [63:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [63:0] _RAND_399;
  reg [63:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [63:0] _RAND_408;
  reg [63:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [63:0] _RAND_417;
  reg [63:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [63:0] _RAND_426;
  reg [63:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [63:0] _RAND_435;
  reg [63:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [63:0] _RAND_444;
  reg [63:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [63:0] _RAND_453;
  reg [63:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [63:0] _RAND_462;
  reg [63:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [63:0] _RAND_471;
  reg [63:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [63:0] _RAND_480;
  reg [63:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [63:0] _RAND_489;
  reg [63:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [63:0] _RAND_498;
  reg [63:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [63:0] _RAND_507;
  reg [63:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [63:0] _RAND_516;
  reg [63:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [63:0] _RAND_525;
  reg [63:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [63:0] _RAND_534;
  reg [63:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [63:0] _RAND_543;
  reg [63:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [63:0] _RAND_552;
  reg [63:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [63:0] _RAND_561;
  reg [63:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [63:0] _RAND_570;
  reg [63:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [63:0] _RAND_579;
  reg [63:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [63:0] _RAND_588;
  reg [63:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [63:0] _RAND_597;
  reg [63:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [63:0] _RAND_606;
  reg [63:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [63:0] _RAND_615;
  reg [63:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [63:0] _RAND_624;
  reg [63:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [63:0] _RAND_633;
  reg [63:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [63:0] _RAND_642;
  reg [63:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
`endif // RANDOMIZE_REG_INIT
  reg [6:0] commit_ptr; // @[rob.scala 46:29]
  reg [6:0] allocate_ptr; // @[rob.scala 47:31]
  reg [1:0] rob_state; // @[rob.scala 53:28]
  reg  last_pc_redirect; // @[rob.scala 55:31]
  wire  _next_rob_state_T_2 = rob_state == 2'h0; // @[rob.scala 215:18]
  wire  _next_rob_state_T_3 = rob_state == 2'h1; // @[rob.scala 216:18]
  wire [6:0] _is_full_T_1 = allocate_ptr + 7'h2; // @[rob.scala 208:30]
  wire [6:0] _is_full_T_4 = allocate_ptr + 7'h1; // @[rob.scala 208:69]
  wire  is_full = _is_full_T_1 == commit_ptr | _is_full_T_4 == commit_ptr; // @[rob.scala 208:52]
  wire  _next_rob_state_T_4 = rob_state == 2'h1 & is_full; // @[rob.scala 216:31]
  wire  _next_rob_state_T_7 = _next_rob_state_T_3 & (io_i_branch_resolve_pack_mispred & io_i_branch_resolve_pack_valid); // @[rob.scala 217:32]
  wire [6:0] _next_rob_state_T_10 = allocate_ptr - 7'h1; // @[rob.scala 218:87]
  wire [7:0] _GEN_41868 = {{1'd0}, _next_rob_state_T_10}; // @[rob.scala 218:71]
  wire [6:0] _next_rob_state_T_13 = allocate_ptr - 7'h2; // @[rob.scala 219:70]
  wire [7:0] _GEN_41869 = {{1'd0}, _next_rob_state_T_13}; // @[rob.scala 219:54]
  wire  _next_rob_state_T_14 = io_i_branch_resolve_pack_rob_idx == _GEN_41869; // @[rob.scala 219:54]
  wire  _next_rob_state_T_16 = rob_state == 2'h2 & (io_i_branch_resolve_pack_rob_idx == _GEN_41868 |
    _next_rob_state_T_14); // @[rob.scala 218:33]
  reg  will_commit_0; // @[rob.scala 89:30]
  wire  _next_rob_state_T_18 = rob_state == 2'h3 & will_commit_0; // @[rob.scala 220:29]
  wire [1:0] _next_rob_state_T_19 = _next_rob_state_T_18 ? 2'h1 : rob_state; // @[Mux.scala 101:16]
  wire [1:0] _next_rob_state_T_20 = _next_rob_state_T_16 ? 2'h1 : _next_rob_state_T_19; // @[Mux.scala 101:16]
  wire [1:0] _next_rob_state_T_21 = _next_rob_state_T_7 ? 2'h2 : _next_rob_state_T_20; // @[Mux.scala 101:16]
  wire [1:0] _next_rob_state_T_22 = _next_rob_state_T_4 ? 2'h3 : _next_rob_state_T_21; // @[Mux.scala 101:16]
  wire [1:0] _next_rob_state_T_23 = _next_rob_state_T_2 ? 2'h1 : _next_rob_state_T_22; // @[Mux.scala 101:16]
  wire [1:0] next_rob_state = io_o_exception | io_i_interrupt | last_pc_redirect ? 2'h0 : _next_rob_state_T_23; // @[rob.scala 214:24]
  wire  _this_num_to_roll_back_T = next_rob_state == 2'h2; // @[rob.scala 74:23]
  wire  _this_num_to_roll_back_T_4 = next_rob_state == 2'h2 & _GEN_41869 > io_i_branch_resolve_pack_rob_idx; // @[rob.scala 74:38]
  wire  _this_num_to_roll_back_T_9 = _this_num_to_roll_back_T & _GEN_41869 == io_i_branch_resolve_pack_rob_idx; // @[rob.scala 75:38]
  wire [1:0] _this_num_to_roll_back_T_17 = _this_num_to_roll_back_T_4 ? 2'h2 : {{1'd0}, _this_num_to_roll_back_T_9}; // @[Mux.scala 101:16]
  reg  rob_valid_0; // @[rob.scala 81:28]
  reg  rob_valid_1; // @[rob.scala 81:28]
  reg  rob_valid_2; // @[rob.scala 81:28]
  reg  rob_valid_3; // @[rob.scala 81:28]
  reg  rob_valid_4; // @[rob.scala 81:28]
  reg  rob_valid_5; // @[rob.scala 81:28]
  reg  rob_valid_6; // @[rob.scala 81:28]
  reg  rob_valid_7; // @[rob.scala 81:28]
  reg  rob_valid_8; // @[rob.scala 81:28]
  reg  rob_valid_9; // @[rob.scala 81:28]
  reg  rob_valid_10; // @[rob.scala 81:28]
  reg  rob_valid_11; // @[rob.scala 81:28]
  reg  rob_valid_12; // @[rob.scala 81:28]
  reg  rob_valid_13; // @[rob.scala 81:28]
  reg  rob_valid_14; // @[rob.scala 81:28]
  reg  rob_valid_15; // @[rob.scala 81:28]
  reg  rob_valid_16; // @[rob.scala 81:28]
  reg  rob_valid_17; // @[rob.scala 81:28]
  reg  rob_valid_18; // @[rob.scala 81:28]
  reg  rob_valid_19; // @[rob.scala 81:28]
  reg  rob_valid_20; // @[rob.scala 81:28]
  reg  rob_valid_21; // @[rob.scala 81:28]
  reg  rob_valid_22; // @[rob.scala 81:28]
  reg  rob_valid_23; // @[rob.scala 81:28]
  reg  rob_valid_24; // @[rob.scala 81:28]
  reg  rob_valid_25; // @[rob.scala 81:28]
  reg  rob_valid_26; // @[rob.scala 81:28]
  reg  rob_valid_27; // @[rob.scala 81:28]
  reg  rob_valid_28; // @[rob.scala 81:28]
  reg  rob_valid_29; // @[rob.scala 81:28]
  reg  rob_valid_30; // @[rob.scala 81:28]
  reg  rob_valid_31; // @[rob.scala 81:28]
  reg  rob_valid_32; // @[rob.scala 81:28]
  reg  rob_valid_33; // @[rob.scala 81:28]
  reg  rob_valid_34; // @[rob.scala 81:28]
  reg  rob_valid_35; // @[rob.scala 81:28]
  reg  rob_valid_36; // @[rob.scala 81:28]
  reg  rob_valid_37; // @[rob.scala 81:28]
  reg  rob_valid_38; // @[rob.scala 81:28]
  reg  rob_valid_39; // @[rob.scala 81:28]
  reg  rob_valid_40; // @[rob.scala 81:28]
  reg  rob_valid_41; // @[rob.scala 81:28]
  reg  rob_valid_42; // @[rob.scala 81:28]
  reg  rob_valid_43; // @[rob.scala 81:28]
  reg  rob_valid_44; // @[rob.scala 81:28]
  reg  rob_valid_45; // @[rob.scala 81:28]
  reg  rob_valid_46; // @[rob.scala 81:28]
  reg  rob_valid_47; // @[rob.scala 81:28]
  reg  rob_valid_48; // @[rob.scala 81:28]
  reg  rob_valid_49; // @[rob.scala 81:28]
  reg  rob_valid_50; // @[rob.scala 81:28]
  reg  rob_valid_51; // @[rob.scala 81:28]
  reg  rob_valid_52; // @[rob.scala 81:28]
  reg  rob_valid_53; // @[rob.scala 81:28]
  reg  rob_valid_54; // @[rob.scala 81:28]
  reg  rob_valid_55; // @[rob.scala 81:28]
  reg  rob_valid_56; // @[rob.scala 81:28]
  reg  rob_valid_57; // @[rob.scala 81:28]
  reg  rob_valid_58; // @[rob.scala 81:28]
  reg  rob_valid_59; // @[rob.scala 81:28]
  reg  rob_valid_60; // @[rob.scala 81:28]
  reg  rob_valid_61; // @[rob.scala 81:28]
  reg  rob_valid_62; // @[rob.scala 81:28]
  reg  rob_valid_63; // @[rob.scala 81:28]
  reg [31:0] rob_uop_0_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_0_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_0_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_0_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_0_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_0_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_0_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_0_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_0_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_1_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_1_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_1_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_1_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_1_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_1_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_1_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_1_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_1_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_2_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_2_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_2_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_2_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_2_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_2_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_2_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_2_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_2_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_3_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_3_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_3_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_3_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_3_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_3_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_3_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_3_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_3_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_4_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_4_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_4_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_4_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_4_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_4_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_4_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_4_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_4_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_5_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_5_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_5_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_5_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_5_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_5_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_5_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_5_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_5_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_6_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_6_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_6_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_6_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_6_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_6_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_6_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_6_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_6_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_7_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_7_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_7_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_7_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_7_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_7_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_7_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_7_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_7_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_8_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_8_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_8_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_8_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_8_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_8_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_8_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_8_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_8_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_9_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_9_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_9_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_9_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_9_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_9_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_9_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_9_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_9_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_10_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_10_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_10_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_10_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_10_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_10_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_10_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_10_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_10_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_11_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_11_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_11_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_11_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_11_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_11_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_11_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_11_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_11_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_12_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_12_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_12_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_12_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_12_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_12_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_12_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_12_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_12_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_13_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_13_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_13_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_13_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_13_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_13_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_13_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_13_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_13_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_14_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_14_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_14_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_14_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_14_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_14_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_14_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_14_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_14_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_15_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_15_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_15_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_15_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_15_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_15_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_15_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_15_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_15_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_16_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_16_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_16_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_16_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_16_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_16_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_16_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_16_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_16_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_17_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_17_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_17_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_17_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_17_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_17_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_17_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_17_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_17_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_18_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_18_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_18_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_18_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_18_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_18_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_18_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_18_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_18_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_19_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_19_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_19_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_19_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_19_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_19_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_19_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_19_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_19_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_20_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_20_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_20_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_20_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_20_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_20_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_20_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_20_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_20_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_21_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_21_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_21_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_21_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_21_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_21_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_21_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_21_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_21_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_22_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_22_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_22_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_22_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_22_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_22_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_22_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_22_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_22_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_23_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_23_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_23_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_23_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_23_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_23_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_23_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_23_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_23_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_24_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_24_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_24_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_24_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_24_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_24_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_24_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_24_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_24_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_25_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_25_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_25_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_25_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_25_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_25_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_25_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_25_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_25_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_26_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_26_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_26_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_26_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_26_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_26_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_26_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_26_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_26_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_27_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_27_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_27_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_27_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_27_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_27_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_27_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_27_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_27_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_28_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_28_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_28_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_28_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_28_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_28_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_28_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_28_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_28_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_29_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_29_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_29_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_29_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_29_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_29_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_29_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_29_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_29_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_30_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_30_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_30_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_30_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_30_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_30_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_30_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_30_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_30_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_31_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_31_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_31_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_31_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_31_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_31_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_31_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_31_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_31_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_32_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_32_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_32_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_32_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_32_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_32_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_32_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_32_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_32_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_33_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_33_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_33_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_33_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_33_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_33_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_33_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_33_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_33_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_34_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_34_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_34_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_34_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_34_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_34_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_34_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_34_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_34_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_35_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_35_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_35_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_35_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_35_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_35_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_35_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_35_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_35_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_36_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_36_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_36_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_36_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_36_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_36_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_36_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_36_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_36_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_37_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_37_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_37_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_37_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_37_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_37_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_37_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_37_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_37_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_38_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_38_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_38_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_38_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_38_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_38_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_38_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_38_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_38_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_39_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_39_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_39_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_39_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_39_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_39_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_39_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_39_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_39_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_40_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_40_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_40_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_40_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_40_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_40_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_40_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_40_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_40_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_41_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_41_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_41_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_41_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_41_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_41_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_41_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_41_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_41_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_42_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_42_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_42_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_42_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_42_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_42_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_42_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_42_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_42_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_43_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_43_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_43_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_43_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_43_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_43_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_43_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_43_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_43_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_44_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_44_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_44_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_44_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_44_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_44_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_44_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_44_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_44_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_45_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_45_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_45_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_45_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_45_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_45_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_45_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_45_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_45_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_46_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_46_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_46_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_46_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_46_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_46_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_46_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_46_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_46_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_47_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_47_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_47_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_47_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_47_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_47_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_47_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_47_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_47_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_48_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_48_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_48_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_48_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_48_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_48_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_48_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_48_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_48_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_49_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_49_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_49_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_49_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_49_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_49_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_49_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_49_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_49_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_50_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_50_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_50_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_50_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_50_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_50_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_50_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_50_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_50_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_51_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_51_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_51_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_51_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_51_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_51_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_51_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_51_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_51_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_52_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_52_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_52_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_52_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_52_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_52_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_52_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_52_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_52_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_53_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_53_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_53_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_53_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_53_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_53_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_53_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_53_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_53_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_54_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_54_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_54_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_54_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_54_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_54_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_54_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_54_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_54_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_55_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_55_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_55_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_55_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_55_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_55_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_55_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_55_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_55_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_56_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_56_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_56_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_56_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_56_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_56_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_56_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_56_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_56_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_57_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_57_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_57_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_57_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_57_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_57_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_57_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_57_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_57_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_58_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_58_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_58_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_58_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_58_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_58_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_58_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_58_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_58_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_59_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_59_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_59_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_59_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_59_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_59_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_59_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_59_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_59_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_60_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_60_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_60_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_60_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_60_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_60_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_60_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_60_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_60_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_61_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_61_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_61_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_61_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_61_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_61_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_61_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_61_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_61_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_62_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_62_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_62_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_62_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_62_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_62_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_62_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_62_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_62_alu_sel; // @[rob.scala 82:26]
  reg [31:0] rob_uop_63_pc; // @[rob.scala 82:26]
  reg [31:0] rob_uop_63_inst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_63_func_code; // @[rob.scala 82:26]
  reg [6:0] rob_uop_63_phy_dst; // @[rob.scala 82:26]
  reg [6:0] rob_uop_63_stale_dst; // @[rob.scala 82:26]
  reg [4:0] rob_uop_63_arch_dst; // @[rob.scala 82:26]
  reg [63:0] rob_uop_63_dst_value; // @[rob.scala 82:26]
  reg [63:0] rob_uop_63_src1_value; // @[rob.scala 82:26]
  reg [4:0] rob_uop_63_alu_sel; // @[rob.scala 82:26]
  reg  rob_done_0; // @[rob.scala 84:27]
  reg  rob_done_1; // @[rob.scala 84:27]
  reg  rob_done_2; // @[rob.scala 84:27]
  reg  rob_done_3; // @[rob.scala 84:27]
  reg  rob_done_4; // @[rob.scala 84:27]
  reg  rob_done_5; // @[rob.scala 84:27]
  reg  rob_done_6; // @[rob.scala 84:27]
  reg  rob_done_7; // @[rob.scala 84:27]
  reg  rob_done_8; // @[rob.scala 84:27]
  reg  rob_done_9; // @[rob.scala 84:27]
  reg  rob_done_10; // @[rob.scala 84:27]
  reg  rob_done_11; // @[rob.scala 84:27]
  reg  rob_done_12; // @[rob.scala 84:27]
  reg  rob_done_13; // @[rob.scala 84:27]
  reg  rob_done_14; // @[rob.scala 84:27]
  reg  rob_done_15; // @[rob.scala 84:27]
  reg  rob_done_16; // @[rob.scala 84:27]
  reg  rob_done_17; // @[rob.scala 84:27]
  reg  rob_done_18; // @[rob.scala 84:27]
  reg  rob_done_19; // @[rob.scala 84:27]
  reg  rob_done_20; // @[rob.scala 84:27]
  reg  rob_done_21; // @[rob.scala 84:27]
  reg  rob_done_22; // @[rob.scala 84:27]
  reg  rob_done_23; // @[rob.scala 84:27]
  reg  rob_done_24; // @[rob.scala 84:27]
  reg  rob_done_25; // @[rob.scala 84:27]
  reg  rob_done_26; // @[rob.scala 84:27]
  reg  rob_done_27; // @[rob.scala 84:27]
  reg  rob_done_28; // @[rob.scala 84:27]
  reg  rob_done_29; // @[rob.scala 84:27]
  reg  rob_done_30; // @[rob.scala 84:27]
  reg  rob_done_31; // @[rob.scala 84:27]
  reg  rob_done_32; // @[rob.scala 84:27]
  reg  rob_done_33; // @[rob.scala 84:27]
  reg  rob_done_34; // @[rob.scala 84:27]
  reg  rob_done_35; // @[rob.scala 84:27]
  reg  rob_done_36; // @[rob.scala 84:27]
  reg  rob_done_37; // @[rob.scala 84:27]
  reg  rob_done_38; // @[rob.scala 84:27]
  reg  rob_done_39; // @[rob.scala 84:27]
  reg  rob_done_40; // @[rob.scala 84:27]
  reg  rob_done_41; // @[rob.scala 84:27]
  reg  rob_done_42; // @[rob.scala 84:27]
  reg  rob_done_43; // @[rob.scala 84:27]
  reg  rob_done_44; // @[rob.scala 84:27]
  reg  rob_done_45; // @[rob.scala 84:27]
  reg  rob_done_46; // @[rob.scala 84:27]
  reg  rob_done_47; // @[rob.scala 84:27]
  reg  rob_done_48; // @[rob.scala 84:27]
  reg  rob_done_49; // @[rob.scala 84:27]
  reg  rob_done_50; // @[rob.scala 84:27]
  reg  rob_done_51; // @[rob.scala 84:27]
  reg  rob_done_52; // @[rob.scala 84:27]
  reg  rob_done_53; // @[rob.scala 84:27]
  reg  rob_done_54; // @[rob.scala 84:27]
  reg  rob_done_55; // @[rob.scala 84:27]
  reg  rob_done_56; // @[rob.scala 84:27]
  reg  rob_done_57; // @[rob.scala 84:27]
  reg  rob_done_58; // @[rob.scala 84:27]
  reg  rob_done_59; // @[rob.scala 84:27]
  reg  rob_done_60; // @[rob.scala 84:27]
  reg  rob_done_61; // @[rob.scala 84:27]
  reg  rob_done_62; // @[rob.scala 84:27]
  reg  rob_done_63; // @[rob.scala 84:27]
  wire  _GEN_1 = 6'h1 == commit_ptr[5:0] ? rob_valid_1 : rob_valid_0; // @[rob.scala 96:{51,51}]
  wire  _GEN_2 = 6'h2 == commit_ptr[5:0] ? rob_valid_2 : _GEN_1; // @[rob.scala 96:{51,51}]
  wire  _GEN_3 = 6'h3 == commit_ptr[5:0] ? rob_valid_3 : _GEN_2; // @[rob.scala 96:{51,51}]
  wire  _GEN_4 = 6'h4 == commit_ptr[5:0] ? rob_valid_4 : _GEN_3; // @[rob.scala 96:{51,51}]
  wire  _GEN_5 = 6'h5 == commit_ptr[5:0] ? rob_valid_5 : _GEN_4; // @[rob.scala 96:{51,51}]
  wire  _GEN_6 = 6'h6 == commit_ptr[5:0] ? rob_valid_6 : _GEN_5; // @[rob.scala 96:{51,51}]
  wire  _GEN_7 = 6'h7 == commit_ptr[5:0] ? rob_valid_7 : _GEN_6; // @[rob.scala 96:{51,51}]
  wire  _GEN_8 = 6'h8 == commit_ptr[5:0] ? rob_valid_8 : _GEN_7; // @[rob.scala 96:{51,51}]
  wire  _GEN_9 = 6'h9 == commit_ptr[5:0] ? rob_valid_9 : _GEN_8; // @[rob.scala 96:{51,51}]
  wire  _GEN_10 = 6'ha == commit_ptr[5:0] ? rob_valid_10 : _GEN_9; // @[rob.scala 96:{51,51}]
  wire  _GEN_11 = 6'hb == commit_ptr[5:0] ? rob_valid_11 : _GEN_10; // @[rob.scala 96:{51,51}]
  wire  _GEN_12 = 6'hc == commit_ptr[5:0] ? rob_valid_12 : _GEN_11; // @[rob.scala 96:{51,51}]
  wire  _GEN_13 = 6'hd == commit_ptr[5:0] ? rob_valid_13 : _GEN_12; // @[rob.scala 96:{51,51}]
  wire  _GEN_14 = 6'he == commit_ptr[5:0] ? rob_valid_14 : _GEN_13; // @[rob.scala 96:{51,51}]
  wire  _GEN_15 = 6'hf == commit_ptr[5:0] ? rob_valid_15 : _GEN_14; // @[rob.scala 96:{51,51}]
  wire  _GEN_16 = 6'h10 == commit_ptr[5:0] ? rob_valid_16 : _GEN_15; // @[rob.scala 96:{51,51}]
  wire  _GEN_17 = 6'h11 == commit_ptr[5:0] ? rob_valid_17 : _GEN_16; // @[rob.scala 96:{51,51}]
  wire  _GEN_18 = 6'h12 == commit_ptr[5:0] ? rob_valid_18 : _GEN_17; // @[rob.scala 96:{51,51}]
  wire  _GEN_19 = 6'h13 == commit_ptr[5:0] ? rob_valid_19 : _GEN_18; // @[rob.scala 96:{51,51}]
  wire  _GEN_20 = 6'h14 == commit_ptr[5:0] ? rob_valid_20 : _GEN_19; // @[rob.scala 96:{51,51}]
  wire  _GEN_21 = 6'h15 == commit_ptr[5:0] ? rob_valid_21 : _GEN_20; // @[rob.scala 96:{51,51}]
  wire  _GEN_22 = 6'h16 == commit_ptr[5:0] ? rob_valid_22 : _GEN_21; // @[rob.scala 96:{51,51}]
  wire  _GEN_23 = 6'h17 == commit_ptr[5:0] ? rob_valid_23 : _GEN_22; // @[rob.scala 96:{51,51}]
  wire  _GEN_24 = 6'h18 == commit_ptr[5:0] ? rob_valid_24 : _GEN_23; // @[rob.scala 96:{51,51}]
  wire  _GEN_25 = 6'h19 == commit_ptr[5:0] ? rob_valid_25 : _GEN_24; // @[rob.scala 96:{51,51}]
  wire  _GEN_26 = 6'h1a == commit_ptr[5:0] ? rob_valid_26 : _GEN_25; // @[rob.scala 96:{51,51}]
  wire  _GEN_27 = 6'h1b == commit_ptr[5:0] ? rob_valid_27 : _GEN_26; // @[rob.scala 96:{51,51}]
  wire  _GEN_28 = 6'h1c == commit_ptr[5:0] ? rob_valid_28 : _GEN_27; // @[rob.scala 96:{51,51}]
  wire  _GEN_29 = 6'h1d == commit_ptr[5:0] ? rob_valid_29 : _GEN_28; // @[rob.scala 96:{51,51}]
  wire  _GEN_30 = 6'h1e == commit_ptr[5:0] ? rob_valid_30 : _GEN_29; // @[rob.scala 96:{51,51}]
  wire  _GEN_31 = 6'h1f == commit_ptr[5:0] ? rob_valid_31 : _GEN_30; // @[rob.scala 96:{51,51}]
  wire  _GEN_32 = 6'h20 == commit_ptr[5:0] ? rob_valid_32 : _GEN_31; // @[rob.scala 96:{51,51}]
  wire  _GEN_33 = 6'h21 == commit_ptr[5:0] ? rob_valid_33 : _GEN_32; // @[rob.scala 96:{51,51}]
  wire  _GEN_34 = 6'h22 == commit_ptr[5:0] ? rob_valid_34 : _GEN_33; // @[rob.scala 96:{51,51}]
  wire  _GEN_35 = 6'h23 == commit_ptr[5:0] ? rob_valid_35 : _GEN_34; // @[rob.scala 96:{51,51}]
  wire  _GEN_36 = 6'h24 == commit_ptr[5:0] ? rob_valid_36 : _GEN_35; // @[rob.scala 96:{51,51}]
  wire  _GEN_37 = 6'h25 == commit_ptr[5:0] ? rob_valid_37 : _GEN_36; // @[rob.scala 96:{51,51}]
  wire  _GEN_38 = 6'h26 == commit_ptr[5:0] ? rob_valid_38 : _GEN_37; // @[rob.scala 96:{51,51}]
  wire  _GEN_39 = 6'h27 == commit_ptr[5:0] ? rob_valid_39 : _GEN_38; // @[rob.scala 96:{51,51}]
  wire  _GEN_40 = 6'h28 == commit_ptr[5:0] ? rob_valid_40 : _GEN_39; // @[rob.scala 96:{51,51}]
  wire  _GEN_41 = 6'h29 == commit_ptr[5:0] ? rob_valid_41 : _GEN_40; // @[rob.scala 96:{51,51}]
  wire  _GEN_42 = 6'h2a == commit_ptr[5:0] ? rob_valid_42 : _GEN_41; // @[rob.scala 96:{51,51}]
  wire  _GEN_43 = 6'h2b == commit_ptr[5:0] ? rob_valid_43 : _GEN_42; // @[rob.scala 96:{51,51}]
  wire  _GEN_44 = 6'h2c == commit_ptr[5:0] ? rob_valid_44 : _GEN_43; // @[rob.scala 96:{51,51}]
  wire  _GEN_45 = 6'h2d == commit_ptr[5:0] ? rob_valid_45 : _GEN_44; // @[rob.scala 96:{51,51}]
  wire  _GEN_46 = 6'h2e == commit_ptr[5:0] ? rob_valid_46 : _GEN_45; // @[rob.scala 96:{51,51}]
  wire  _GEN_47 = 6'h2f == commit_ptr[5:0] ? rob_valid_47 : _GEN_46; // @[rob.scala 96:{51,51}]
  wire  _GEN_48 = 6'h30 == commit_ptr[5:0] ? rob_valid_48 : _GEN_47; // @[rob.scala 96:{51,51}]
  wire  _GEN_49 = 6'h31 == commit_ptr[5:0] ? rob_valid_49 : _GEN_48; // @[rob.scala 96:{51,51}]
  wire  _GEN_50 = 6'h32 == commit_ptr[5:0] ? rob_valid_50 : _GEN_49; // @[rob.scala 96:{51,51}]
  wire  _GEN_51 = 6'h33 == commit_ptr[5:0] ? rob_valid_51 : _GEN_50; // @[rob.scala 96:{51,51}]
  wire  _GEN_52 = 6'h34 == commit_ptr[5:0] ? rob_valid_52 : _GEN_51; // @[rob.scala 96:{51,51}]
  wire  _GEN_53 = 6'h35 == commit_ptr[5:0] ? rob_valid_53 : _GEN_52; // @[rob.scala 96:{51,51}]
  wire  _GEN_54 = 6'h36 == commit_ptr[5:0] ? rob_valid_54 : _GEN_53; // @[rob.scala 96:{51,51}]
  wire  _GEN_55 = 6'h37 == commit_ptr[5:0] ? rob_valid_55 : _GEN_54; // @[rob.scala 96:{51,51}]
  wire  _GEN_56 = 6'h38 == commit_ptr[5:0] ? rob_valid_56 : _GEN_55; // @[rob.scala 96:{51,51}]
  wire  _GEN_57 = 6'h39 == commit_ptr[5:0] ? rob_valid_57 : _GEN_56; // @[rob.scala 96:{51,51}]
  wire  _GEN_58 = 6'h3a == commit_ptr[5:0] ? rob_valid_58 : _GEN_57; // @[rob.scala 96:{51,51}]
  wire  _GEN_59 = 6'h3b == commit_ptr[5:0] ? rob_valid_59 : _GEN_58; // @[rob.scala 96:{51,51}]
  wire  _GEN_60 = 6'h3c == commit_ptr[5:0] ? rob_valid_60 : _GEN_59; // @[rob.scala 96:{51,51}]
  wire  _GEN_61 = 6'h3d == commit_ptr[5:0] ? rob_valid_61 : _GEN_60; // @[rob.scala 96:{51,51}]
  wire  _GEN_62 = 6'h3e == commit_ptr[5:0] ? rob_valid_62 : _GEN_61; // @[rob.scala 96:{51,51}]
  wire  _GEN_63 = 6'h3f == commit_ptr[5:0] ? rob_valid_63 : _GEN_62; // @[rob.scala 96:{51,51}]
  wire  _GEN_65 = 6'h1 == commit_ptr[5:0] ? rob_done_1 : rob_done_0; // @[rob.scala 96:{51,51}]
  wire  _GEN_66 = 6'h2 == commit_ptr[5:0] ? rob_done_2 : _GEN_65; // @[rob.scala 96:{51,51}]
  wire  _GEN_67 = 6'h3 == commit_ptr[5:0] ? rob_done_3 : _GEN_66; // @[rob.scala 96:{51,51}]
  wire  _GEN_68 = 6'h4 == commit_ptr[5:0] ? rob_done_4 : _GEN_67; // @[rob.scala 96:{51,51}]
  wire  _GEN_69 = 6'h5 == commit_ptr[5:0] ? rob_done_5 : _GEN_68; // @[rob.scala 96:{51,51}]
  wire  _GEN_70 = 6'h6 == commit_ptr[5:0] ? rob_done_6 : _GEN_69; // @[rob.scala 96:{51,51}]
  wire  _GEN_71 = 6'h7 == commit_ptr[5:0] ? rob_done_7 : _GEN_70; // @[rob.scala 96:{51,51}]
  wire  _GEN_72 = 6'h8 == commit_ptr[5:0] ? rob_done_8 : _GEN_71; // @[rob.scala 96:{51,51}]
  wire  _GEN_73 = 6'h9 == commit_ptr[5:0] ? rob_done_9 : _GEN_72; // @[rob.scala 96:{51,51}]
  wire  _GEN_74 = 6'ha == commit_ptr[5:0] ? rob_done_10 : _GEN_73; // @[rob.scala 96:{51,51}]
  wire  _GEN_75 = 6'hb == commit_ptr[5:0] ? rob_done_11 : _GEN_74; // @[rob.scala 96:{51,51}]
  wire  _GEN_76 = 6'hc == commit_ptr[5:0] ? rob_done_12 : _GEN_75; // @[rob.scala 96:{51,51}]
  wire  _GEN_77 = 6'hd == commit_ptr[5:0] ? rob_done_13 : _GEN_76; // @[rob.scala 96:{51,51}]
  wire  _GEN_78 = 6'he == commit_ptr[5:0] ? rob_done_14 : _GEN_77; // @[rob.scala 96:{51,51}]
  wire  _GEN_79 = 6'hf == commit_ptr[5:0] ? rob_done_15 : _GEN_78; // @[rob.scala 96:{51,51}]
  wire  _GEN_80 = 6'h10 == commit_ptr[5:0] ? rob_done_16 : _GEN_79; // @[rob.scala 96:{51,51}]
  wire  _GEN_81 = 6'h11 == commit_ptr[5:0] ? rob_done_17 : _GEN_80; // @[rob.scala 96:{51,51}]
  wire  _GEN_82 = 6'h12 == commit_ptr[5:0] ? rob_done_18 : _GEN_81; // @[rob.scala 96:{51,51}]
  wire  _GEN_83 = 6'h13 == commit_ptr[5:0] ? rob_done_19 : _GEN_82; // @[rob.scala 96:{51,51}]
  wire  _GEN_84 = 6'h14 == commit_ptr[5:0] ? rob_done_20 : _GEN_83; // @[rob.scala 96:{51,51}]
  wire  _GEN_85 = 6'h15 == commit_ptr[5:0] ? rob_done_21 : _GEN_84; // @[rob.scala 96:{51,51}]
  wire  _GEN_86 = 6'h16 == commit_ptr[5:0] ? rob_done_22 : _GEN_85; // @[rob.scala 96:{51,51}]
  wire  _GEN_87 = 6'h17 == commit_ptr[5:0] ? rob_done_23 : _GEN_86; // @[rob.scala 96:{51,51}]
  wire  _GEN_88 = 6'h18 == commit_ptr[5:0] ? rob_done_24 : _GEN_87; // @[rob.scala 96:{51,51}]
  wire  _GEN_89 = 6'h19 == commit_ptr[5:0] ? rob_done_25 : _GEN_88; // @[rob.scala 96:{51,51}]
  wire  _GEN_90 = 6'h1a == commit_ptr[5:0] ? rob_done_26 : _GEN_89; // @[rob.scala 96:{51,51}]
  wire  _GEN_91 = 6'h1b == commit_ptr[5:0] ? rob_done_27 : _GEN_90; // @[rob.scala 96:{51,51}]
  wire  _GEN_92 = 6'h1c == commit_ptr[5:0] ? rob_done_28 : _GEN_91; // @[rob.scala 96:{51,51}]
  wire  _GEN_93 = 6'h1d == commit_ptr[5:0] ? rob_done_29 : _GEN_92; // @[rob.scala 96:{51,51}]
  wire  _GEN_94 = 6'h1e == commit_ptr[5:0] ? rob_done_30 : _GEN_93; // @[rob.scala 96:{51,51}]
  wire  _GEN_95 = 6'h1f == commit_ptr[5:0] ? rob_done_31 : _GEN_94; // @[rob.scala 96:{51,51}]
  wire  _GEN_96 = 6'h20 == commit_ptr[5:0] ? rob_done_32 : _GEN_95; // @[rob.scala 96:{51,51}]
  wire  _GEN_97 = 6'h21 == commit_ptr[5:0] ? rob_done_33 : _GEN_96; // @[rob.scala 96:{51,51}]
  wire  _GEN_98 = 6'h22 == commit_ptr[5:0] ? rob_done_34 : _GEN_97; // @[rob.scala 96:{51,51}]
  wire  _GEN_99 = 6'h23 == commit_ptr[5:0] ? rob_done_35 : _GEN_98; // @[rob.scala 96:{51,51}]
  wire  _GEN_100 = 6'h24 == commit_ptr[5:0] ? rob_done_36 : _GEN_99; // @[rob.scala 96:{51,51}]
  wire  _GEN_101 = 6'h25 == commit_ptr[5:0] ? rob_done_37 : _GEN_100; // @[rob.scala 96:{51,51}]
  wire  _GEN_102 = 6'h26 == commit_ptr[5:0] ? rob_done_38 : _GEN_101; // @[rob.scala 96:{51,51}]
  wire  _GEN_103 = 6'h27 == commit_ptr[5:0] ? rob_done_39 : _GEN_102; // @[rob.scala 96:{51,51}]
  wire  _GEN_104 = 6'h28 == commit_ptr[5:0] ? rob_done_40 : _GEN_103; // @[rob.scala 96:{51,51}]
  wire  _GEN_105 = 6'h29 == commit_ptr[5:0] ? rob_done_41 : _GEN_104; // @[rob.scala 96:{51,51}]
  wire  _GEN_106 = 6'h2a == commit_ptr[5:0] ? rob_done_42 : _GEN_105; // @[rob.scala 96:{51,51}]
  wire  _GEN_107 = 6'h2b == commit_ptr[5:0] ? rob_done_43 : _GEN_106; // @[rob.scala 96:{51,51}]
  wire  _GEN_108 = 6'h2c == commit_ptr[5:0] ? rob_done_44 : _GEN_107; // @[rob.scala 96:{51,51}]
  wire  _GEN_109 = 6'h2d == commit_ptr[5:0] ? rob_done_45 : _GEN_108; // @[rob.scala 96:{51,51}]
  wire  _GEN_110 = 6'h2e == commit_ptr[5:0] ? rob_done_46 : _GEN_109; // @[rob.scala 96:{51,51}]
  wire  _GEN_111 = 6'h2f == commit_ptr[5:0] ? rob_done_47 : _GEN_110; // @[rob.scala 96:{51,51}]
  wire  _GEN_112 = 6'h30 == commit_ptr[5:0] ? rob_done_48 : _GEN_111; // @[rob.scala 96:{51,51}]
  wire  _GEN_113 = 6'h31 == commit_ptr[5:0] ? rob_done_49 : _GEN_112; // @[rob.scala 96:{51,51}]
  wire  _GEN_114 = 6'h32 == commit_ptr[5:0] ? rob_done_50 : _GEN_113; // @[rob.scala 96:{51,51}]
  wire  _GEN_115 = 6'h33 == commit_ptr[5:0] ? rob_done_51 : _GEN_114; // @[rob.scala 96:{51,51}]
  wire  _GEN_116 = 6'h34 == commit_ptr[5:0] ? rob_done_52 : _GEN_115; // @[rob.scala 96:{51,51}]
  wire  _GEN_117 = 6'h35 == commit_ptr[5:0] ? rob_done_53 : _GEN_116; // @[rob.scala 96:{51,51}]
  wire  _GEN_118 = 6'h36 == commit_ptr[5:0] ? rob_done_54 : _GEN_117; // @[rob.scala 96:{51,51}]
  wire  _GEN_119 = 6'h37 == commit_ptr[5:0] ? rob_done_55 : _GEN_118; // @[rob.scala 96:{51,51}]
  wire  _GEN_120 = 6'h38 == commit_ptr[5:0] ? rob_done_56 : _GEN_119; // @[rob.scala 96:{51,51}]
  wire  _GEN_121 = 6'h39 == commit_ptr[5:0] ? rob_done_57 : _GEN_120; // @[rob.scala 96:{51,51}]
  wire  _GEN_122 = 6'h3a == commit_ptr[5:0] ? rob_done_58 : _GEN_121; // @[rob.scala 96:{51,51}]
  wire  _GEN_123 = 6'h3b == commit_ptr[5:0] ? rob_done_59 : _GEN_122; // @[rob.scala 96:{51,51}]
  wire  _GEN_124 = 6'h3c == commit_ptr[5:0] ? rob_done_60 : _GEN_123; // @[rob.scala 96:{51,51}]
  wire  _GEN_125 = 6'h3d == commit_ptr[5:0] ? rob_done_61 : _GEN_124; // @[rob.scala 96:{51,51}]
  wire  _GEN_126 = 6'h3e == commit_ptr[5:0] ? rob_done_62 : _GEN_125; // @[rob.scala 96:{51,51}]
  wire  _GEN_127 = 6'h3f == commit_ptr[5:0] ? rob_done_63 : _GEN_126; // @[rob.scala 96:{51,51}]
  wire  next_can_commit_0 = _GEN_63 & _GEN_127; // @[rob.scala 96:51]
  wire [6:0] _next_can_commit_1_T_1 = commit_ptr + 7'h1; // @[rob.scala 97:47]
  wire  _GEN_129 = 6'h1 == _next_can_commit_1_T_1[5:0] ? rob_valid_1 : rob_valid_0; // @[rob.scala 97:{53,53}]
  wire  _GEN_130 = 6'h2 == _next_can_commit_1_T_1[5:0] ? rob_valid_2 : _GEN_129; // @[rob.scala 97:{53,53}]
  wire  _GEN_131 = 6'h3 == _next_can_commit_1_T_1[5:0] ? rob_valid_3 : _GEN_130; // @[rob.scala 97:{53,53}]
  wire  _GEN_132 = 6'h4 == _next_can_commit_1_T_1[5:0] ? rob_valid_4 : _GEN_131; // @[rob.scala 97:{53,53}]
  wire  _GEN_133 = 6'h5 == _next_can_commit_1_T_1[5:0] ? rob_valid_5 : _GEN_132; // @[rob.scala 97:{53,53}]
  wire  _GEN_134 = 6'h6 == _next_can_commit_1_T_1[5:0] ? rob_valid_6 : _GEN_133; // @[rob.scala 97:{53,53}]
  wire  _GEN_135 = 6'h7 == _next_can_commit_1_T_1[5:0] ? rob_valid_7 : _GEN_134; // @[rob.scala 97:{53,53}]
  wire  _GEN_136 = 6'h8 == _next_can_commit_1_T_1[5:0] ? rob_valid_8 : _GEN_135; // @[rob.scala 97:{53,53}]
  wire  _GEN_137 = 6'h9 == _next_can_commit_1_T_1[5:0] ? rob_valid_9 : _GEN_136; // @[rob.scala 97:{53,53}]
  wire  _GEN_138 = 6'ha == _next_can_commit_1_T_1[5:0] ? rob_valid_10 : _GEN_137; // @[rob.scala 97:{53,53}]
  wire  _GEN_139 = 6'hb == _next_can_commit_1_T_1[5:0] ? rob_valid_11 : _GEN_138; // @[rob.scala 97:{53,53}]
  wire  _GEN_140 = 6'hc == _next_can_commit_1_T_1[5:0] ? rob_valid_12 : _GEN_139; // @[rob.scala 97:{53,53}]
  wire  _GEN_141 = 6'hd == _next_can_commit_1_T_1[5:0] ? rob_valid_13 : _GEN_140; // @[rob.scala 97:{53,53}]
  wire  _GEN_142 = 6'he == _next_can_commit_1_T_1[5:0] ? rob_valid_14 : _GEN_141; // @[rob.scala 97:{53,53}]
  wire  _GEN_143 = 6'hf == _next_can_commit_1_T_1[5:0] ? rob_valid_15 : _GEN_142; // @[rob.scala 97:{53,53}]
  wire  _GEN_144 = 6'h10 == _next_can_commit_1_T_1[5:0] ? rob_valid_16 : _GEN_143; // @[rob.scala 97:{53,53}]
  wire  _GEN_145 = 6'h11 == _next_can_commit_1_T_1[5:0] ? rob_valid_17 : _GEN_144; // @[rob.scala 97:{53,53}]
  wire  _GEN_146 = 6'h12 == _next_can_commit_1_T_1[5:0] ? rob_valid_18 : _GEN_145; // @[rob.scala 97:{53,53}]
  wire  _GEN_147 = 6'h13 == _next_can_commit_1_T_1[5:0] ? rob_valid_19 : _GEN_146; // @[rob.scala 97:{53,53}]
  wire  _GEN_148 = 6'h14 == _next_can_commit_1_T_1[5:0] ? rob_valid_20 : _GEN_147; // @[rob.scala 97:{53,53}]
  wire  _GEN_149 = 6'h15 == _next_can_commit_1_T_1[5:0] ? rob_valid_21 : _GEN_148; // @[rob.scala 97:{53,53}]
  wire  _GEN_150 = 6'h16 == _next_can_commit_1_T_1[5:0] ? rob_valid_22 : _GEN_149; // @[rob.scala 97:{53,53}]
  wire  _GEN_151 = 6'h17 == _next_can_commit_1_T_1[5:0] ? rob_valid_23 : _GEN_150; // @[rob.scala 97:{53,53}]
  wire  _GEN_152 = 6'h18 == _next_can_commit_1_T_1[5:0] ? rob_valid_24 : _GEN_151; // @[rob.scala 97:{53,53}]
  wire  _GEN_153 = 6'h19 == _next_can_commit_1_T_1[5:0] ? rob_valid_25 : _GEN_152; // @[rob.scala 97:{53,53}]
  wire  _GEN_154 = 6'h1a == _next_can_commit_1_T_1[5:0] ? rob_valid_26 : _GEN_153; // @[rob.scala 97:{53,53}]
  wire  _GEN_155 = 6'h1b == _next_can_commit_1_T_1[5:0] ? rob_valid_27 : _GEN_154; // @[rob.scala 97:{53,53}]
  wire  _GEN_156 = 6'h1c == _next_can_commit_1_T_1[5:0] ? rob_valid_28 : _GEN_155; // @[rob.scala 97:{53,53}]
  wire  _GEN_157 = 6'h1d == _next_can_commit_1_T_1[5:0] ? rob_valid_29 : _GEN_156; // @[rob.scala 97:{53,53}]
  wire  _GEN_158 = 6'h1e == _next_can_commit_1_T_1[5:0] ? rob_valid_30 : _GEN_157; // @[rob.scala 97:{53,53}]
  wire  _GEN_159 = 6'h1f == _next_can_commit_1_T_1[5:0] ? rob_valid_31 : _GEN_158; // @[rob.scala 97:{53,53}]
  wire  _GEN_160 = 6'h20 == _next_can_commit_1_T_1[5:0] ? rob_valid_32 : _GEN_159; // @[rob.scala 97:{53,53}]
  wire  _GEN_161 = 6'h21 == _next_can_commit_1_T_1[5:0] ? rob_valid_33 : _GEN_160; // @[rob.scala 97:{53,53}]
  wire  _GEN_162 = 6'h22 == _next_can_commit_1_T_1[5:0] ? rob_valid_34 : _GEN_161; // @[rob.scala 97:{53,53}]
  wire  _GEN_163 = 6'h23 == _next_can_commit_1_T_1[5:0] ? rob_valid_35 : _GEN_162; // @[rob.scala 97:{53,53}]
  wire  _GEN_164 = 6'h24 == _next_can_commit_1_T_1[5:0] ? rob_valid_36 : _GEN_163; // @[rob.scala 97:{53,53}]
  wire  _GEN_165 = 6'h25 == _next_can_commit_1_T_1[5:0] ? rob_valid_37 : _GEN_164; // @[rob.scala 97:{53,53}]
  wire  _GEN_166 = 6'h26 == _next_can_commit_1_T_1[5:0] ? rob_valid_38 : _GEN_165; // @[rob.scala 97:{53,53}]
  wire  _GEN_167 = 6'h27 == _next_can_commit_1_T_1[5:0] ? rob_valid_39 : _GEN_166; // @[rob.scala 97:{53,53}]
  wire  _GEN_168 = 6'h28 == _next_can_commit_1_T_1[5:0] ? rob_valid_40 : _GEN_167; // @[rob.scala 97:{53,53}]
  wire  _GEN_169 = 6'h29 == _next_can_commit_1_T_1[5:0] ? rob_valid_41 : _GEN_168; // @[rob.scala 97:{53,53}]
  wire  _GEN_170 = 6'h2a == _next_can_commit_1_T_1[5:0] ? rob_valid_42 : _GEN_169; // @[rob.scala 97:{53,53}]
  wire  _GEN_171 = 6'h2b == _next_can_commit_1_T_1[5:0] ? rob_valid_43 : _GEN_170; // @[rob.scala 97:{53,53}]
  wire  _GEN_172 = 6'h2c == _next_can_commit_1_T_1[5:0] ? rob_valid_44 : _GEN_171; // @[rob.scala 97:{53,53}]
  wire  _GEN_173 = 6'h2d == _next_can_commit_1_T_1[5:0] ? rob_valid_45 : _GEN_172; // @[rob.scala 97:{53,53}]
  wire  _GEN_174 = 6'h2e == _next_can_commit_1_T_1[5:0] ? rob_valid_46 : _GEN_173; // @[rob.scala 97:{53,53}]
  wire  _GEN_175 = 6'h2f == _next_can_commit_1_T_1[5:0] ? rob_valid_47 : _GEN_174; // @[rob.scala 97:{53,53}]
  wire  _GEN_176 = 6'h30 == _next_can_commit_1_T_1[5:0] ? rob_valid_48 : _GEN_175; // @[rob.scala 97:{53,53}]
  wire  _GEN_177 = 6'h31 == _next_can_commit_1_T_1[5:0] ? rob_valid_49 : _GEN_176; // @[rob.scala 97:{53,53}]
  wire  _GEN_178 = 6'h32 == _next_can_commit_1_T_1[5:0] ? rob_valid_50 : _GEN_177; // @[rob.scala 97:{53,53}]
  wire  _GEN_179 = 6'h33 == _next_can_commit_1_T_1[5:0] ? rob_valid_51 : _GEN_178; // @[rob.scala 97:{53,53}]
  wire  _GEN_180 = 6'h34 == _next_can_commit_1_T_1[5:0] ? rob_valid_52 : _GEN_179; // @[rob.scala 97:{53,53}]
  wire  _GEN_181 = 6'h35 == _next_can_commit_1_T_1[5:0] ? rob_valid_53 : _GEN_180; // @[rob.scala 97:{53,53}]
  wire  _GEN_182 = 6'h36 == _next_can_commit_1_T_1[5:0] ? rob_valid_54 : _GEN_181; // @[rob.scala 97:{53,53}]
  wire  _GEN_183 = 6'h37 == _next_can_commit_1_T_1[5:0] ? rob_valid_55 : _GEN_182; // @[rob.scala 97:{53,53}]
  wire  _GEN_184 = 6'h38 == _next_can_commit_1_T_1[5:0] ? rob_valid_56 : _GEN_183; // @[rob.scala 97:{53,53}]
  wire  _GEN_185 = 6'h39 == _next_can_commit_1_T_1[5:0] ? rob_valid_57 : _GEN_184; // @[rob.scala 97:{53,53}]
  wire  _GEN_186 = 6'h3a == _next_can_commit_1_T_1[5:0] ? rob_valid_58 : _GEN_185; // @[rob.scala 97:{53,53}]
  wire  _GEN_187 = 6'h3b == _next_can_commit_1_T_1[5:0] ? rob_valid_59 : _GEN_186; // @[rob.scala 97:{53,53}]
  wire  _GEN_188 = 6'h3c == _next_can_commit_1_T_1[5:0] ? rob_valid_60 : _GEN_187; // @[rob.scala 97:{53,53}]
  wire  _GEN_189 = 6'h3d == _next_can_commit_1_T_1[5:0] ? rob_valid_61 : _GEN_188; // @[rob.scala 97:{53,53}]
  wire  _GEN_190 = 6'h3e == _next_can_commit_1_T_1[5:0] ? rob_valid_62 : _GEN_189; // @[rob.scala 97:{53,53}]
  wire  _GEN_191 = 6'h3f == _next_can_commit_1_T_1[5:0] ? rob_valid_63 : _GEN_190; // @[rob.scala 97:{53,53}]
  wire  _GEN_193 = 6'h1 == _next_can_commit_1_T_1[5:0] ? rob_done_1 : rob_done_0; // @[rob.scala 97:{53,53}]
  wire  _GEN_194 = 6'h2 == _next_can_commit_1_T_1[5:0] ? rob_done_2 : _GEN_193; // @[rob.scala 97:{53,53}]
  wire  _GEN_195 = 6'h3 == _next_can_commit_1_T_1[5:0] ? rob_done_3 : _GEN_194; // @[rob.scala 97:{53,53}]
  wire  _GEN_196 = 6'h4 == _next_can_commit_1_T_1[5:0] ? rob_done_4 : _GEN_195; // @[rob.scala 97:{53,53}]
  wire  _GEN_197 = 6'h5 == _next_can_commit_1_T_1[5:0] ? rob_done_5 : _GEN_196; // @[rob.scala 97:{53,53}]
  wire  _GEN_198 = 6'h6 == _next_can_commit_1_T_1[5:0] ? rob_done_6 : _GEN_197; // @[rob.scala 97:{53,53}]
  wire  _GEN_199 = 6'h7 == _next_can_commit_1_T_1[5:0] ? rob_done_7 : _GEN_198; // @[rob.scala 97:{53,53}]
  wire  _GEN_200 = 6'h8 == _next_can_commit_1_T_1[5:0] ? rob_done_8 : _GEN_199; // @[rob.scala 97:{53,53}]
  wire  _GEN_201 = 6'h9 == _next_can_commit_1_T_1[5:0] ? rob_done_9 : _GEN_200; // @[rob.scala 97:{53,53}]
  wire  _GEN_202 = 6'ha == _next_can_commit_1_T_1[5:0] ? rob_done_10 : _GEN_201; // @[rob.scala 97:{53,53}]
  wire  _GEN_203 = 6'hb == _next_can_commit_1_T_1[5:0] ? rob_done_11 : _GEN_202; // @[rob.scala 97:{53,53}]
  wire  _GEN_204 = 6'hc == _next_can_commit_1_T_1[5:0] ? rob_done_12 : _GEN_203; // @[rob.scala 97:{53,53}]
  wire  _GEN_205 = 6'hd == _next_can_commit_1_T_1[5:0] ? rob_done_13 : _GEN_204; // @[rob.scala 97:{53,53}]
  wire  _GEN_206 = 6'he == _next_can_commit_1_T_1[5:0] ? rob_done_14 : _GEN_205; // @[rob.scala 97:{53,53}]
  wire  _GEN_207 = 6'hf == _next_can_commit_1_T_1[5:0] ? rob_done_15 : _GEN_206; // @[rob.scala 97:{53,53}]
  wire  _GEN_208 = 6'h10 == _next_can_commit_1_T_1[5:0] ? rob_done_16 : _GEN_207; // @[rob.scala 97:{53,53}]
  wire  _GEN_209 = 6'h11 == _next_can_commit_1_T_1[5:0] ? rob_done_17 : _GEN_208; // @[rob.scala 97:{53,53}]
  wire  _GEN_210 = 6'h12 == _next_can_commit_1_T_1[5:0] ? rob_done_18 : _GEN_209; // @[rob.scala 97:{53,53}]
  wire  _GEN_211 = 6'h13 == _next_can_commit_1_T_1[5:0] ? rob_done_19 : _GEN_210; // @[rob.scala 97:{53,53}]
  wire  _GEN_212 = 6'h14 == _next_can_commit_1_T_1[5:0] ? rob_done_20 : _GEN_211; // @[rob.scala 97:{53,53}]
  wire  _GEN_213 = 6'h15 == _next_can_commit_1_T_1[5:0] ? rob_done_21 : _GEN_212; // @[rob.scala 97:{53,53}]
  wire  _GEN_214 = 6'h16 == _next_can_commit_1_T_1[5:0] ? rob_done_22 : _GEN_213; // @[rob.scala 97:{53,53}]
  wire  _GEN_215 = 6'h17 == _next_can_commit_1_T_1[5:0] ? rob_done_23 : _GEN_214; // @[rob.scala 97:{53,53}]
  wire  _GEN_216 = 6'h18 == _next_can_commit_1_T_1[5:0] ? rob_done_24 : _GEN_215; // @[rob.scala 97:{53,53}]
  wire  _GEN_217 = 6'h19 == _next_can_commit_1_T_1[5:0] ? rob_done_25 : _GEN_216; // @[rob.scala 97:{53,53}]
  wire  _GEN_218 = 6'h1a == _next_can_commit_1_T_1[5:0] ? rob_done_26 : _GEN_217; // @[rob.scala 97:{53,53}]
  wire  _GEN_219 = 6'h1b == _next_can_commit_1_T_1[5:0] ? rob_done_27 : _GEN_218; // @[rob.scala 97:{53,53}]
  wire  _GEN_220 = 6'h1c == _next_can_commit_1_T_1[5:0] ? rob_done_28 : _GEN_219; // @[rob.scala 97:{53,53}]
  wire  _GEN_221 = 6'h1d == _next_can_commit_1_T_1[5:0] ? rob_done_29 : _GEN_220; // @[rob.scala 97:{53,53}]
  wire  _GEN_222 = 6'h1e == _next_can_commit_1_T_1[5:0] ? rob_done_30 : _GEN_221; // @[rob.scala 97:{53,53}]
  wire  _GEN_223 = 6'h1f == _next_can_commit_1_T_1[5:0] ? rob_done_31 : _GEN_222; // @[rob.scala 97:{53,53}]
  wire  _GEN_224 = 6'h20 == _next_can_commit_1_T_1[5:0] ? rob_done_32 : _GEN_223; // @[rob.scala 97:{53,53}]
  wire  _GEN_225 = 6'h21 == _next_can_commit_1_T_1[5:0] ? rob_done_33 : _GEN_224; // @[rob.scala 97:{53,53}]
  wire  _GEN_226 = 6'h22 == _next_can_commit_1_T_1[5:0] ? rob_done_34 : _GEN_225; // @[rob.scala 97:{53,53}]
  wire  _GEN_227 = 6'h23 == _next_can_commit_1_T_1[5:0] ? rob_done_35 : _GEN_226; // @[rob.scala 97:{53,53}]
  wire  _GEN_228 = 6'h24 == _next_can_commit_1_T_1[5:0] ? rob_done_36 : _GEN_227; // @[rob.scala 97:{53,53}]
  wire  _GEN_229 = 6'h25 == _next_can_commit_1_T_1[5:0] ? rob_done_37 : _GEN_228; // @[rob.scala 97:{53,53}]
  wire  _GEN_230 = 6'h26 == _next_can_commit_1_T_1[5:0] ? rob_done_38 : _GEN_229; // @[rob.scala 97:{53,53}]
  wire  _GEN_231 = 6'h27 == _next_can_commit_1_T_1[5:0] ? rob_done_39 : _GEN_230; // @[rob.scala 97:{53,53}]
  wire  _GEN_232 = 6'h28 == _next_can_commit_1_T_1[5:0] ? rob_done_40 : _GEN_231; // @[rob.scala 97:{53,53}]
  wire  _GEN_233 = 6'h29 == _next_can_commit_1_T_1[5:0] ? rob_done_41 : _GEN_232; // @[rob.scala 97:{53,53}]
  wire  _GEN_234 = 6'h2a == _next_can_commit_1_T_1[5:0] ? rob_done_42 : _GEN_233; // @[rob.scala 97:{53,53}]
  wire  _GEN_235 = 6'h2b == _next_can_commit_1_T_1[5:0] ? rob_done_43 : _GEN_234; // @[rob.scala 97:{53,53}]
  wire  _GEN_236 = 6'h2c == _next_can_commit_1_T_1[5:0] ? rob_done_44 : _GEN_235; // @[rob.scala 97:{53,53}]
  wire  _GEN_237 = 6'h2d == _next_can_commit_1_T_1[5:0] ? rob_done_45 : _GEN_236; // @[rob.scala 97:{53,53}]
  wire  _GEN_238 = 6'h2e == _next_can_commit_1_T_1[5:0] ? rob_done_46 : _GEN_237; // @[rob.scala 97:{53,53}]
  wire  _GEN_239 = 6'h2f == _next_can_commit_1_T_1[5:0] ? rob_done_47 : _GEN_238; // @[rob.scala 97:{53,53}]
  wire  _GEN_240 = 6'h30 == _next_can_commit_1_T_1[5:0] ? rob_done_48 : _GEN_239; // @[rob.scala 97:{53,53}]
  wire  _GEN_241 = 6'h31 == _next_can_commit_1_T_1[5:0] ? rob_done_49 : _GEN_240; // @[rob.scala 97:{53,53}]
  wire  _GEN_242 = 6'h32 == _next_can_commit_1_T_1[5:0] ? rob_done_50 : _GEN_241; // @[rob.scala 97:{53,53}]
  wire  _GEN_243 = 6'h33 == _next_can_commit_1_T_1[5:0] ? rob_done_51 : _GEN_242; // @[rob.scala 97:{53,53}]
  wire  _GEN_244 = 6'h34 == _next_can_commit_1_T_1[5:0] ? rob_done_52 : _GEN_243; // @[rob.scala 97:{53,53}]
  wire  _GEN_245 = 6'h35 == _next_can_commit_1_T_1[5:0] ? rob_done_53 : _GEN_244; // @[rob.scala 97:{53,53}]
  wire  _GEN_246 = 6'h36 == _next_can_commit_1_T_1[5:0] ? rob_done_54 : _GEN_245; // @[rob.scala 97:{53,53}]
  wire  _GEN_247 = 6'h37 == _next_can_commit_1_T_1[5:0] ? rob_done_55 : _GEN_246; // @[rob.scala 97:{53,53}]
  wire  _GEN_248 = 6'h38 == _next_can_commit_1_T_1[5:0] ? rob_done_56 : _GEN_247; // @[rob.scala 97:{53,53}]
  wire  _GEN_249 = 6'h39 == _next_can_commit_1_T_1[5:0] ? rob_done_57 : _GEN_248; // @[rob.scala 97:{53,53}]
  wire  _GEN_250 = 6'h3a == _next_can_commit_1_T_1[5:0] ? rob_done_58 : _GEN_249; // @[rob.scala 97:{53,53}]
  wire  _GEN_251 = 6'h3b == _next_can_commit_1_T_1[5:0] ? rob_done_59 : _GEN_250; // @[rob.scala 97:{53,53}]
  wire  _GEN_252 = 6'h3c == _next_can_commit_1_T_1[5:0] ? rob_done_60 : _GEN_251; // @[rob.scala 97:{53,53}]
  wire  _GEN_253 = 6'h3d == _next_can_commit_1_T_1[5:0] ? rob_done_61 : _GEN_252; // @[rob.scala 97:{53,53}]
  wire  _GEN_254 = 6'h3e == _next_can_commit_1_T_1[5:0] ? rob_done_62 : _GEN_253; // @[rob.scala 97:{53,53}]
  wire  _GEN_255 = 6'h3f == _next_can_commit_1_T_1[5:0] ? rob_done_63 : _GEN_254; // @[rob.scala 97:{53,53}]
  wire  next_can_commit_1 = _GEN_191 & _GEN_255; // @[rob.scala 97:53]
  wire  _next_will_commit_0_T = ~io_i_interrupt; // @[rob.scala 99:28]
  wire  _next_will_commit_0_T_5 = next_rob_state == 2'h1; // @[rob.scala 99:114]
  wire  _next_will_commit_0_T_6 = next_rob_state == 2'h3; // @[rob.scala 99:143]
  wire  _next_will_commit_0_T_7 = next_rob_state == 2'h1 | next_rob_state == 2'h3; // @[rob.scala 99:126]
  wire  next_will_commit_0 = ~io_i_interrupt & next_can_commit_0 & (next_rob_state == 2'h1 | next_rob_state == 2'h3); // @[rob.scala 99:96]
  wire [6:0] _GEN_321 = 6'h1 == commit_ptr[5:0] ? rob_uop_1_func_code : rob_uop_0_func_code; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_322 = 6'h2 == commit_ptr[5:0] ? rob_uop_2_func_code : _GEN_321; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_323 = 6'h3 == commit_ptr[5:0] ? rob_uop_3_func_code : _GEN_322; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_324 = 6'h4 == commit_ptr[5:0] ? rob_uop_4_func_code : _GEN_323; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_325 = 6'h5 == commit_ptr[5:0] ? rob_uop_5_func_code : _GEN_324; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_326 = 6'h6 == commit_ptr[5:0] ? rob_uop_6_func_code : _GEN_325; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_327 = 6'h7 == commit_ptr[5:0] ? rob_uop_7_func_code : _GEN_326; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_328 = 6'h8 == commit_ptr[5:0] ? rob_uop_8_func_code : _GEN_327; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_329 = 6'h9 == commit_ptr[5:0] ? rob_uop_9_func_code : _GEN_328; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_330 = 6'ha == commit_ptr[5:0] ? rob_uop_10_func_code : _GEN_329; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_331 = 6'hb == commit_ptr[5:0] ? rob_uop_11_func_code : _GEN_330; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_332 = 6'hc == commit_ptr[5:0] ? rob_uop_12_func_code : _GEN_331; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_333 = 6'hd == commit_ptr[5:0] ? rob_uop_13_func_code : _GEN_332; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_334 = 6'he == commit_ptr[5:0] ? rob_uop_14_func_code : _GEN_333; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_335 = 6'hf == commit_ptr[5:0] ? rob_uop_15_func_code : _GEN_334; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_336 = 6'h10 == commit_ptr[5:0] ? rob_uop_16_func_code : _GEN_335; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_337 = 6'h11 == commit_ptr[5:0] ? rob_uop_17_func_code : _GEN_336; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_338 = 6'h12 == commit_ptr[5:0] ? rob_uop_18_func_code : _GEN_337; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_339 = 6'h13 == commit_ptr[5:0] ? rob_uop_19_func_code : _GEN_338; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_340 = 6'h14 == commit_ptr[5:0] ? rob_uop_20_func_code : _GEN_339; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_341 = 6'h15 == commit_ptr[5:0] ? rob_uop_21_func_code : _GEN_340; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_342 = 6'h16 == commit_ptr[5:0] ? rob_uop_22_func_code : _GEN_341; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_343 = 6'h17 == commit_ptr[5:0] ? rob_uop_23_func_code : _GEN_342; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_344 = 6'h18 == commit_ptr[5:0] ? rob_uop_24_func_code : _GEN_343; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_345 = 6'h19 == commit_ptr[5:0] ? rob_uop_25_func_code : _GEN_344; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_346 = 6'h1a == commit_ptr[5:0] ? rob_uop_26_func_code : _GEN_345; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_347 = 6'h1b == commit_ptr[5:0] ? rob_uop_27_func_code : _GEN_346; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_348 = 6'h1c == commit_ptr[5:0] ? rob_uop_28_func_code : _GEN_347; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_349 = 6'h1d == commit_ptr[5:0] ? rob_uop_29_func_code : _GEN_348; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_350 = 6'h1e == commit_ptr[5:0] ? rob_uop_30_func_code : _GEN_349; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_351 = 6'h1f == commit_ptr[5:0] ? rob_uop_31_func_code : _GEN_350; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_352 = 6'h20 == commit_ptr[5:0] ? rob_uop_32_func_code : _GEN_351; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_353 = 6'h21 == commit_ptr[5:0] ? rob_uop_33_func_code : _GEN_352; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_354 = 6'h22 == commit_ptr[5:0] ? rob_uop_34_func_code : _GEN_353; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_355 = 6'h23 == commit_ptr[5:0] ? rob_uop_35_func_code : _GEN_354; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_356 = 6'h24 == commit_ptr[5:0] ? rob_uop_36_func_code : _GEN_355; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_357 = 6'h25 == commit_ptr[5:0] ? rob_uop_37_func_code : _GEN_356; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_358 = 6'h26 == commit_ptr[5:0] ? rob_uop_38_func_code : _GEN_357; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_359 = 6'h27 == commit_ptr[5:0] ? rob_uop_39_func_code : _GEN_358; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_360 = 6'h28 == commit_ptr[5:0] ? rob_uop_40_func_code : _GEN_359; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_361 = 6'h29 == commit_ptr[5:0] ? rob_uop_41_func_code : _GEN_360; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_362 = 6'h2a == commit_ptr[5:0] ? rob_uop_42_func_code : _GEN_361; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_363 = 6'h2b == commit_ptr[5:0] ? rob_uop_43_func_code : _GEN_362; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_364 = 6'h2c == commit_ptr[5:0] ? rob_uop_44_func_code : _GEN_363; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_365 = 6'h2d == commit_ptr[5:0] ? rob_uop_45_func_code : _GEN_364; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_366 = 6'h2e == commit_ptr[5:0] ? rob_uop_46_func_code : _GEN_365; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_367 = 6'h2f == commit_ptr[5:0] ? rob_uop_47_func_code : _GEN_366; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_368 = 6'h30 == commit_ptr[5:0] ? rob_uop_48_func_code : _GEN_367; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_369 = 6'h31 == commit_ptr[5:0] ? rob_uop_49_func_code : _GEN_368; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_370 = 6'h32 == commit_ptr[5:0] ? rob_uop_50_func_code : _GEN_369; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_371 = 6'h33 == commit_ptr[5:0] ? rob_uop_51_func_code : _GEN_370; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_372 = 6'h34 == commit_ptr[5:0] ? rob_uop_52_func_code : _GEN_371; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_373 = 6'h35 == commit_ptr[5:0] ? rob_uop_53_func_code : _GEN_372; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_374 = 6'h36 == commit_ptr[5:0] ? rob_uop_54_func_code : _GEN_373; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_375 = 6'h37 == commit_ptr[5:0] ? rob_uop_55_func_code : _GEN_374; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_376 = 6'h38 == commit_ptr[5:0] ? rob_uop_56_func_code : _GEN_375; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_377 = 6'h39 == commit_ptr[5:0] ? rob_uop_57_func_code : _GEN_376; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_378 = 6'h3a == commit_ptr[5:0] ? rob_uop_58_func_code : _GEN_377; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_379 = 6'h3b == commit_ptr[5:0] ? rob_uop_59_func_code : _GEN_378; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_380 = 6'h3c == commit_ptr[5:0] ? rob_uop_60_func_code : _GEN_379; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_381 = 6'h3d == commit_ptr[5:0] ? rob_uop_61_func_code : _GEN_380; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_382 = 6'h3e == commit_ptr[5:0] ? rob_uop_62_func_code : _GEN_381; // @[rob.scala 100:{79,79}]
  wire [6:0] _GEN_383 = 6'h3f == commit_ptr[5:0] ? rob_uop_63_func_code : _GEN_382; // @[rob.scala 100:{79,79}]
  wire [4:0] _GEN_385 = 6'h1 == commit_ptr[5:0] ? rob_uop_1_alu_sel : rob_uop_0_alu_sel; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_386 = 6'h2 == commit_ptr[5:0] ? rob_uop_2_alu_sel : _GEN_385; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_387 = 6'h3 == commit_ptr[5:0] ? rob_uop_3_alu_sel : _GEN_386; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_388 = 6'h4 == commit_ptr[5:0] ? rob_uop_4_alu_sel : _GEN_387; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_389 = 6'h5 == commit_ptr[5:0] ? rob_uop_5_alu_sel : _GEN_388; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_390 = 6'h6 == commit_ptr[5:0] ? rob_uop_6_alu_sel : _GEN_389; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_391 = 6'h7 == commit_ptr[5:0] ? rob_uop_7_alu_sel : _GEN_390; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_392 = 6'h8 == commit_ptr[5:0] ? rob_uop_8_alu_sel : _GEN_391; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_393 = 6'h9 == commit_ptr[5:0] ? rob_uop_9_alu_sel : _GEN_392; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_394 = 6'ha == commit_ptr[5:0] ? rob_uop_10_alu_sel : _GEN_393; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_395 = 6'hb == commit_ptr[5:0] ? rob_uop_11_alu_sel : _GEN_394; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_396 = 6'hc == commit_ptr[5:0] ? rob_uop_12_alu_sel : _GEN_395; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_397 = 6'hd == commit_ptr[5:0] ? rob_uop_13_alu_sel : _GEN_396; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_398 = 6'he == commit_ptr[5:0] ? rob_uop_14_alu_sel : _GEN_397; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_399 = 6'hf == commit_ptr[5:0] ? rob_uop_15_alu_sel : _GEN_398; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_400 = 6'h10 == commit_ptr[5:0] ? rob_uop_16_alu_sel : _GEN_399; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_401 = 6'h11 == commit_ptr[5:0] ? rob_uop_17_alu_sel : _GEN_400; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_402 = 6'h12 == commit_ptr[5:0] ? rob_uop_18_alu_sel : _GEN_401; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_403 = 6'h13 == commit_ptr[5:0] ? rob_uop_19_alu_sel : _GEN_402; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_404 = 6'h14 == commit_ptr[5:0] ? rob_uop_20_alu_sel : _GEN_403; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_405 = 6'h15 == commit_ptr[5:0] ? rob_uop_21_alu_sel : _GEN_404; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_406 = 6'h16 == commit_ptr[5:0] ? rob_uop_22_alu_sel : _GEN_405; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_407 = 6'h17 == commit_ptr[5:0] ? rob_uop_23_alu_sel : _GEN_406; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_408 = 6'h18 == commit_ptr[5:0] ? rob_uop_24_alu_sel : _GEN_407; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_409 = 6'h19 == commit_ptr[5:0] ? rob_uop_25_alu_sel : _GEN_408; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_410 = 6'h1a == commit_ptr[5:0] ? rob_uop_26_alu_sel : _GEN_409; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_411 = 6'h1b == commit_ptr[5:0] ? rob_uop_27_alu_sel : _GEN_410; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_412 = 6'h1c == commit_ptr[5:0] ? rob_uop_28_alu_sel : _GEN_411; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_413 = 6'h1d == commit_ptr[5:0] ? rob_uop_29_alu_sel : _GEN_412; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_414 = 6'h1e == commit_ptr[5:0] ? rob_uop_30_alu_sel : _GEN_413; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_415 = 6'h1f == commit_ptr[5:0] ? rob_uop_31_alu_sel : _GEN_414; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_416 = 6'h20 == commit_ptr[5:0] ? rob_uop_32_alu_sel : _GEN_415; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_417 = 6'h21 == commit_ptr[5:0] ? rob_uop_33_alu_sel : _GEN_416; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_418 = 6'h22 == commit_ptr[5:0] ? rob_uop_34_alu_sel : _GEN_417; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_419 = 6'h23 == commit_ptr[5:0] ? rob_uop_35_alu_sel : _GEN_418; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_420 = 6'h24 == commit_ptr[5:0] ? rob_uop_36_alu_sel : _GEN_419; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_421 = 6'h25 == commit_ptr[5:0] ? rob_uop_37_alu_sel : _GEN_420; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_422 = 6'h26 == commit_ptr[5:0] ? rob_uop_38_alu_sel : _GEN_421; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_423 = 6'h27 == commit_ptr[5:0] ? rob_uop_39_alu_sel : _GEN_422; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_424 = 6'h28 == commit_ptr[5:0] ? rob_uop_40_alu_sel : _GEN_423; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_425 = 6'h29 == commit_ptr[5:0] ? rob_uop_41_alu_sel : _GEN_424; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_426 = 6'h2a == commit_ptr[5:0] ? rob_uop_42_alu_sel : _GEN_425; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_427 = 6'h2b == commit_ptr[5:0] ? rob_uop_43_alu_sel : _GEN_426; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_428 = 6'h2c == commit_ptr[5:0] ? rob_uop_44_alu_sel : _GEN_427; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_429 = 6'h2d == commit_ptr[5:0] ? rob_uop_45_alu_sel : _GEN_428; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_430 = 6'h2e == commit_ptr[5:0] ? rob_uop_46_alu_sel : _GEN_429; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_431 = 6'h2f == commit_ptr[5:0] ? rob_uop_47_alu_sel : _GEN_430; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_432 = 6'h30 == commit_ptr[5:0] ? rob_uop_48_alu_sel : _GEN_431; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_433 = 6'h31 == commit_ptr[5:0] ? rob_uop_49_alu_sel : _GEN_432; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_434 = 6'h32 == commit_ptr[5:0] ? rob_uop_50_alu_sel : _GEN_433; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_435 = 6'h33 == commit_ptr[5:0] ? rob_uop_51_alu_sel : _GEN_434; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_436 = 6'h34 == commit_ptr[5:0] ? rob_uop_52_alu_sel : _GEN_435; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_437 = 6'h35 == commit_ptr[5:0] ? rob_uop_53_alu_sel : _GEN_436; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_438 = 6'h36 == commit_ptr[5:0] ? rob_uop_54_alu_sel : _GEN_437; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_439 = 6'h37 == commit_ptr[5:0] ? rob_uop_55_alu_sel : _GEN_438; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_440 = 6'h38 == commit_ptr[5:0] ? rob_uop_56_alu_sel : _GEN_439; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_441 = 6'h39 == commit_ptr[5:0] ? rob_uop_57_alu_sel : _GEN_440; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_442 = 6'h3a == commit_ptr[5:0] ? rob_uop_58_alu_sel : _GEN_441; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_443 = 6'h3b == commit_ptr[5:0] ? rob_uop_59_alu_sel : _GEN_442; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_444 = 6'h3c == commit_ptr[5:0] ? rob_uop_60_alu_sel : _GEN_443; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_445 = 6'h3d == commit_ptr[5:0] ? rob_uop_61_alu_sel : _GEN_444; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_446 = 6'h3e == commit_ptr[5:0] ? rob_uop_62_alu_sel : _GEN_445; // @[rob.scala 101:{39,39}]
  wire [4:0] _GEN_447 = 6'h3f == commit_ptr[5:0] ? rob_uop_63_alu_sel : _GEN_446; // @[rob.scala 101:{39,39}]
  wire  _next_will_commit_1_T_10 = _GEN_447 == 5'h4 | _GEN_447 == 5'h6 | _GEN_447 == 5'h5; // @[rob.scala 101:102]
  wire  _next_will_commit_1_T_13 = _next_will_commit_0_T & ~(_GEN_383 == 7'h20 & _next_will_commit_1_T_10); // @[rob.scala 100:44]
  wire  next_will_commit_1 = _next_will_commit_1_T_13 & next_can_commit_0 & next_can_commit_1 & _next_will_commit_0_T_7; // @[rob.scala 102:114]
  wire [31:0] _GEN_769 = 6'h1 == commit_ptr[5:0] ? rob_uop_1_pc : rob_uop_0_pc; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_770 = 6'h2 == commit_ptr[5:0] ? rob_uop_2_pc : _GEN_769; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_771 = 6'h3 == commit_ptr[5:0] ? rob_uop_3_pc : _GEN_770; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_772 = 6'h4 == commit_ptr[5:0] ? rob_uop_4_pc : _GEN_771; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_773 = 6'h5 == commit_ptr[5:0] ? rob_uop_5_pc : _GEN_772; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_774 = 6'h6 == commit_ptr[5:0] ? rob_uop_6_pc : _GEN_773; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_775 = 6'h7 == commit_ptr[5:0] ? rob_uop_7_pc : _GEN_774; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_776 = 6'h8 == commit_ptr[5:0] ? rob_uop_8_pc : _GEN_775; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_777 = 6'h9 == commit_ptr[5:0] ? rob_uop_9_pc : _GEN_776; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_778 = 6'ha == commit_ptr[5:0] ? rob_uop_10_pc : _GEN_777; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_779 = 6'hb == commit_ptr[5:0] ? rob_uop_11_pc : _GEN_778; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_780 = 6'hc == commit_ptr[5:0] ? rob_uop_12_pc : _GEN_779; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_781 = 6'hd == commit_ptr[5:0] ? rob_uop_13_pc : _GEN_780; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_782 = 6'he == commit_ptr[5:0] ? rob_uop_14_pc : _GEN_781; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_783 = 6'hf == commit_ptr[5:0] ? rob_uop_15_pc : _GEN_782; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_784 = 6'h10 == commit_ptr[5:0] ? rob_uop_16_pc : _GEN_783; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_785 = 6'h11 == commit_ptr[5:0] ? rob_uop_17_pc : _GEN_784; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_786 = 6'h12 == commit_ptr[5:0] ? rob_uop_18_pc : _GEN_785; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_787 = 6'h13 == commit_ptr[5:0] ? rob_uop_19_pc : _GEN_786; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_788 = 6'h14 == commit_ptr[5:0] ? rob_uop_20_pc : _GEN_787; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_789 = 6'h15 == commit_ptr[5:0] ? rob_uop_21_pc : _GEN_788; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_790 = 6'h16 == commit_ptr[5:0] ? rob_uop_22_pc : _GEN_789; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_791 = 6'h17 == commit_ptr[5:0] ? rob_uop_23_pc : _GEN_790; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_792 = 6'h18 == commit_ptr[5:0] ? rob_uop_24_pc : _GEN_791; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_793 = 6'h19 == commit_ptr[5:0] ? rob_uop_25_pc : _GEN_792; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_794 = 6'h1a == commit_ptr[5:0] ? rob_uop_26_pc : _GEN_793; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_795 = 6'h1b == commit_ptr[5:0] ? rob_uop_27_pc : _GEN_794; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_796 = 6'h1c == commit_ptr[5:0] ? rob_uop_28_pc : _GEN_795; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_797 = 6'h1d == commit_ptr[5:0] ? rob_uop_29_pc : _GEN_796; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_798 = 6'h1e == commit_ptr[5:0] ? rob_uop_30_pc : _GEN_797; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_799 = 6'h1f == commit_ptr[5:0] ? rob_uop_31_pc : _GEN_798; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_800 = 6'h20 == commit_ptr[5:0] ? rob_uop_32_pc : _GEN_799; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_801 = 6'h21 == commit_ptr[5:0] ? rob_uop_33_pc : _GEN_800; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_802 = 6'h22 == commit_ptr[5:0] ? rob_uop_34_pc : _GEN_801; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_803 = 6'h23 == commit_ptr[5:0] ? rob_uop_35_pc : _GEN_802; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_804 = 6'h24 == commit_ptr[5:0] ? rob_uop_36_pc : _GEN_803; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_805 = 6'h25 == commit_ptr[5:0] ? rob_uop_37_pc : _GEN_804; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_806 = 6'h26 == commit_ptr[5:0] ? rob_uop_38_pc : _GEN_805; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_807 = 6'h27 == commit_ptr[5:0] ? rob_uop_39_pc : _GEN_806; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_808 = 6'h28 == commit_ptr[5:0] ? rob_uop_40_pc : _GEN_807; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_809 = 6'h29 == commit_ptr[5:0] ? rob_uop_41_pc : _GEN_808; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_810 = 6'h2a == commit_ptr[5:0] ? rob_uop_42_pc : _GEN_809; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_811 = 6'h2b == commit_ptr[5:0] ? rob_uop_43_pc : _GEN_810; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_812 = 6'h2c == commit_ptr[5:0] ? rob_uop_44_pc : _GEN_811; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_813 = 6'h2d == commit_ptr[5:0] ? rob_uop_45_pc : _GEN_812; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_814 = 6'h2e == commit_ptr[5:0] ? rob_uop_46_pc : _GEN_813; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_815 = 6'h2f == commit_ptr[5:0] ? rob_uop_47_pc : _GEN_814; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_816 = 6'h30 == commit_ptr[5:0] ? rob_uop_48_pc : _GEN_815; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_817 = 6'h31 == commit_ptr[5:0] ? rob_uop_49_pc : _GEN_816; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_818 = 6'h32 == commit_ptr[5:0] ? rob_uop_50_pc : _GEN_817; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_819 = 6'h33 == commit_ptr[5:0] ? rob_uop_51_pc : _GEN_818; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_820 = 6'h34 == commit_ptr[5:0] ? rob_uop_52_pc : _GEN_819; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_821 = 6'h35 == commit_ptr[5:0] ? rob_uop_53_pc : _GEN_820; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_822 = 6'h36 == commit_ptr[5:0] ? rob_uop_54_pc : _GEN_821; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_823 = 6'h37 == commit_ptr[5:0] ? rob_uop_55_pc : _GEN_822; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_824 = 6'h38 == commit_ptr[5:0] ? rob_uop_56_pc : _GEN_823; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_825 = 6'h39 == commit_ptr[5:0] ? rob_uop_57_pc : _GEN_824; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_826 = 6'h3a == commit_ptr[5:0] ? rob_uop_58_pc : _GEN_825; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_827 = 6'h3b == commit_ptr[5:0] ? rob_uop_59_pc : _GEN_826; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_828 = 6'h3c == commit_ptr[5:0] ? rob_uop_60_pc : _GEN_827; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_829 = 6'h3d == commit_ptr[5:0] ? rob_uop_61_pc : _GEN_828; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_830 = 6'h3e == commit_ptr[5:0] ? rob_uop_62_pc : _GEN_829; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_833 = 6'h1 == commit_ptr[5:0] ? rob_uop_1_inst : rob_uop_0_inst; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_834 = 6'h2 == commit_ptr[5:0] ? rob_uop_2_inst : _GEN_833; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_835 = 6'h3 == commit_ptr[5:0] ? rob_uop_3_inst : _GEN_834; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_836 = 6'h4 == commit_ptr[5:0] ? rob_uop_4_inst : _GEN_835; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_837 = 6'h5 == commit_ptr[5:0] ? rob_uop_5_inst : _GEN_836; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_838 = 6'h6 == commit_ptr[5:0] ? rob_uop_6_inst : _GEN_837; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_839 = 6'h7 == commit_ptr[5:0] ? rob_uop_7_inst : _GEN_838; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_840 = 6'h8 == commit_ptr[5:0] ? rob_uop_8_inst : _GEN_839; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_841 = 6'h9 == commit_ptr[5:0] ? rob_uop_9_inst : _GEN_840; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_842 = 6'ha == commit_ptr[5:0] ? rob_uop_10_inst : _GEN_841; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_843 = 6'hb == commit_ptr[5:0] ? rob_uop_11_inst : _GEN_842; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_844 = 6'hc == commit_ptr[5:0] ? rob_uop_12_inst : _GEN_843; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_845 = 6'hd == commit_ptr[5:0] ? rob_uop_13_inst : _GEN_844; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_846 = 6'he == commit_ptr[5:0] ? rob_uop_14_inst : _GEN_845; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_847 = 6'hf == commit_ptr[5:0] ? rob_uop_15_inst : _GEN_846; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_848 = 6'h10 == commit_ptr[5:0] ? rob_uop_16_inst : _GEN_847; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_849 = 6'h11 == commit_ptr[5:0] ? rob_uop_17_inst : _GEN_848; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_850 = 6'h12 == commit_ptr[5:0] ? rob_uop_18_inst : _GEN_849; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_851 = 6'h13 == commit_ptr[5:0] ? rob_uop_19_inst : _GEN_850; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_852 = 6'h14 == commit_ptr[5:0] ? rob_uop_20_inst : _GEN_851; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_853 = 6'h15 == commit_ptr[5:0] ? rob_uop_21_inst : _GEN_852; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_854 = 6'h16 == commit_ptr[5:0] ? rob_uop_22_inst : _GEN_853; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_855 = 6'h17 == commit_ptr[5:0] ? rob_uop_23_inst : _GEN_854; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_856 = 6'h18 == commit_ptr[5:0] ? rob_uop_24_inst : _GEN_855; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_857 = 6'h19 == commit_ptr[5:0] ? rob_uop_25_inst : _GEN_856; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_858 = 6'h1a == commit_ptr[5:0] ? rob_uop_26_inst : _GEN_857; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_859 = 6'h1b == commit_ptr[5:0] ? rob_uop_27_inst : _GEN_858; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_860 = 6'h1c == commit_ptr[5:0] ? rob_uop_28_inst : _GEN_859; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_861 = 6'h1d == commit_ptr[5:0] ? rob_uop_29_inst : _GEN_860; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_862 = 6'h1e == commit_ptr[5:0] ? rob_uop_30_inst : _GEN_861; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_863 = 6'h1f == commit_ptr[5:0] ? rob_uop_31_inst : _GEN_862; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_864 = 6'h20 == commit_ptr[5:0] ? rob_uop_32_inst : _GEN_863; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_865 = 6'h21 == commit_ptr[5:0] ? rob_uop_33_inst : _GEN_864; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_866 = 6'h22 == commit_ptr[5:0] ? rob_uop_34_inst : _GEN_865; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_867 = 6'h23 == commit_ptr[5:0] ? rob_uop_35_inst : _GEN_866; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_868 = 6'h24 == commit_ptr[5:0] ? rob_uop_36_inst : _GEN_867; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_869 = 6'h25 == commit_ptr[5:0] ? rob_uop_37_inst : _GEN_868; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_870 = 6'h26 == commit_ptr[5:0] ? rob_uop_38_inst : _GEN_869; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_871 = 6'h27 == commit_ptr[5:0] ? rob_uop_39_inst : _GEN_870; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_872 = 6'h28 == commit_ptr[5:0] ? rob_uop_40_inst : _GEN_871; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_873 = 6'h29 == commit_ptr[5:0] ? rob_uop_41_inst : _GEN_872; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_874 = 6'h2a == commit_ptr[5:0] ? rob_uop_42_inst : _GEN_873; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_875 = 6'h2b == commit_ptr[5:0] ? rob_uop_43_inst : _GEN_874; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_876 = 6'h2c == commit_ptr[5:0] ? rob_uop_44_inst : _GEN_875; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_877 = 6'h2d == commit_ptr[5:0] ? rob_uop_45_inst : _GEN_876; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_878 = 6'h2e == commit_ptr[5:0] ? rob_uop_46_inst : _GEN_877; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_879 = 6'h2f == commit_ptr[5:0] ? rob_uop_47_inst : _GEN_878; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_880 = 6'h30 == commit_ptr[5:0] ? rob_uop_48_inst : _GEN_879; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_881 = 6'h31 == commit_ptr[5:0] ? rob_uop_49_inst : _GEN_880; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_882 = 6'h32 == commit_ptr[5:0] ? rob_uop_50_inst : _GEN_881; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_883 = 6'h33 == commit_ptr[5:0] ? rob_uop_51_inst : _GEN_882; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_884 = 6'h34 == commit_ptr[5:0] ? rob_uop_52_inst : _GEN_883; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_885 = 6'h35 == commit_ptr[5:0] ? rob_uop_53_inst : _GEN_884; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_886 = 6'h36 == commit_ptr[5:0] ? rob_uop_54_inst : _GEN_885; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_887 = 6'h37 == commit_ptr[5:0] ? rob_uop_55_inst : _GEN_886; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_888 = 6'h38 == commit_ptr[5:0] ? rob_uop_56_inst : _GEN_887; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_889 = 6'h39 == commit_ptr[5:0] ? rob_uop_57_inst : _GEN_888; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_890 = 6'h3a == commit_ptr[5:0] ? rob_uop_58_inst : _GEN_889; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_891 = 6'h3b == commit_ptr[5:0] ? rob_uop_59_inst : _GEN_890; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_892 = 6'h3c == commit_ptr[5:0] ? rob_uop_60_inst : _GEN_891; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_893 = 6'h3d == commit_ptr[5:0] ? rob_uop_61_inst : _GEN_892; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_894 = 6'h3e == commit_ptr[5:0] ? rob_uop_62_inst : _GEN_893; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1281 = 6'h1 == commit_ptr[5:0] ? rob_uop_1_phy_dst : rob_uop_0_phy_dst; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1282 = 6'h2 == commit_ptr[5:0] ? rob_uop_2_phy_dst : _GEN_1281; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1283 = 6'h3 == commit_ptr[5:0] ? rob_uop_3_phy_dst : _GEN_1282; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1284 = 6'h4 == commit_ptr[5:0] ? rob_uop_4_phy_dst : _GEN_1283; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1285 = 6'h5 == commit_ptr[5:0] ? rob_uop_5_phy_dst : _GEN_1284; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1286 = 6'h6 == commit_ptr[5:0] ? rob_uop_6_phy_dst : _GEN_1285; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1287 = 6'h7 == commit_ptr[5:0] ? rob_uop_7_phy_dst : _GEN_1286; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1288 = 6'h8 == commit_ptr[5:0] ? rob_uop_8_phy_dst : _GEN_1287; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1289 = 6'h9 == commit_ptr[5:0] ? rob_uop_9_phy_dst : _GEN_1288; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1290 = 6'ha == commit_ptr[5:0] ? rob_uop_10_phy_dst : _GEN_1289; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1291 = 6'hb == commit_ptr[5:0] ? rob_uop_11_phy_dst : _GEN_1290; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1292 = 6'hc == commit_ptr[5:0] ? rob_uop_12_phy_dst : _GEN_1291; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1293 = 6'hd == commit_ptr[5:0] ? rob_uop_13_phy_dst : _GEN_1292; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1294 = 6'he == commit_ptr[5:0] ? rob_uop_14_phy_dst : _GEN_1293; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1295 = 6'hf == commit_ptr[5:0] ? rob_uop_15_phy_dst : _GEN_1294; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1296 = 6'h10 == commit_ptr[5:0] ? rob_uop_16_phy_dst : _GEN_1295; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1297 = 6'h11 == commit_ptr[5:0] ? rob_uop_17_phy_dst : _GEN_1296; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1298 = 6'h12 == commit_ptr[5:0] ? rob_uop_18_phy_dst : _GEN_1297; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1299 = 6'h13 == commit_ptr[5:0] ? rob_uop_19_phy_dst : _GEN_1298; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1300 = 6'h14 == commit_ptr[5:0] ? rob_uop_20_phy_dst : _GEN_1299; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1301 = 6'h15 == commit_ptr[5:0] ? rob_uop_21_phy_dst : _GEN_1300; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1302 = 6'h16 == commit_ptr[5:0] ? rob_uop_22_phy_dst : _GEN_1301; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1303 = 6'h17 == commit_ptr[5:0] ? rob_uop_23_phy_dst : _GEN_1302; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1304 = 6'h18 == commit_ptr[5:0] ? rob_uop_24_phy_dst : _GEN_1303; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1305 = 6'h19 == commit_ptr[5:0] ? rob_uop_25_phy_dst : _GEN_1304; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1306 = 6'h1a == commit_ptr[5:0] ? rob_uop_26_phy_dst : _GEN_1305; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1307 = 6'h1b == commit_ptr[5:0] ? rob_uop_27_phy_dst : _GEN_1306; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1308 = 6'h1c == commit_ptr[5:0] ? rob_uop_28_phy_dst : _GEN_1307; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1309 = 6'h1d == commit_ptr[5:0] ? rob_uop_29_phy_dst : _GEN_1308; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1310 = 6'h1e == commit_ptr[5:0] ? rob_uop_30_phy_dst : _GEN_1309; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1311 = 6'h1f == commit_ptr[5:0] ? rob_uop_31_phy_dst : _GEN_1310; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1312 = 6'h20 == commit_ptr[5:0] ? rob_uop_32_phy_dst : _GEN_1311; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1313 = 6'h21 == commit_ptr[5:0] ? rob_uop_33_phy_dst : _GEN_1312; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1314 = 6'h22 == commit_ptr[5:0] ? rob_uop_34_phy_dst : _GEN_1313; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1315 = 6'h23 == commit_ptr[5:0] ? rob_uop_35_phy_dst : _GEN_1314; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1316 = 6'h24 == commit_ptr[5:0] ? rob_uop_36_phy_dst : _GEN_1315; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1317 = 6'h25 == commit_ptr[5:0] ? rob_uop_37_phy_dst : _GEN_1316; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1318 = 6'h26 == commit_ptr[5:0] ? rob_uop_38_phy_dst : _GEN_1317; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1319 = 6'h27 == commit_ptr[5:0] ? rob_uop_39_phy_dst : _GEN_1318; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1320 = 6'h28 == commit_ptr[5:0] ? rob_uop_40_phy_dst : _GEN_1319; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1321 = 6'h29 == commit_ptr[5:0] ? rob_uop_41_phy_dst : _GEN_1320; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1322 = 6'h2a == commit_ptr[5:0] ? rob_uop_42_phy_dst : _GEN_1321; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1323 = 6'h2b == commit_ptr[5:0] ? rob_uop_43_phy_dst : _GEN_1322; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1324 = 6'h2c == commit_ptr[5:0] ? rob_uop_44_phy_dst : _GEN_1323; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1325 = 6'h2d == commit_ptr[5:0] ? rob_uop_45_phy_dst : _GEN_1324; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1326 = 6'h2e == commit_ptr[5:0] ? rob_uop_46_phy_dst : _GEN_1325; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1327 = 6'h2f == commit_ptr[5:0] ? rob_uop_47_phy_dst : _GEN_1326; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1328 = 6'h30 == commit_ptr[5:0] ? rob_uop_48_phy_dst : _GEN_1327; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1329 = 6'h31 == commit_ptr[5:0] ? rob_uop_49_phy_dst : _GEN_1328; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1330 = 6'h32 == commit_ptr[5:0] ? rob_uop_50_phy_dst : _GEN_1329; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1331 = 6'h33 == commit_ptr[5:0] ? rob_uop_51_phy_dst : _GEN_1330; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1332 = 6'h34 == commit_ptr[5:0] ? rob_uop_52_phy_dst : _GEN_1331; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1333 = 6'h35 == commit_ptr[5:0] ? rob_uop_53_phy_dst : _GEN_1332; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1334 = 6'h36 == commit_ptr[5:0] ? rob_uop_54_phy_dst : _GEN_1333; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1335 = 6'h37 == commit_ptr[5:0] ? rob_uop_55_phy_dst : _GEN_1334; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1336 = 6'h38 == commit_ptr[5:0] ? rob_uop_56_phy_dst : _GEN_1335; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1337 = 6'h39 == commit_ptr[5:0] ? rob_uop_57_phy_dst : _GEN_1336; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1338 = 6'h3a == commit_ptr[5:0] ? rob_uop_58_phy_dst : _GEN_1337; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1339 = 6'h3b == commit_ptr[5:0] ? rob_uop_59_phy_dst : _GEN_1338; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1340 = 6'h3c == commit_ptr[5:0] ? rob_uop_60_phy_dst : _GEN_1339; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1341 = 6'h3d == commit_ptr[5:0] ? rob_uop_61_phy_dst : _GEN_1340; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1342 = 6'h3e == commit_ptr[5:0] ? rob_uop_62_phy_dst : _GEN_1341; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1345 = 6'h1 == commit_ptr[5:0] ? rob_uop_1_stale_dst : rob_uop_0_stale_dst; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1346 = 6'h2 == commit_ptr[5:0] ? rob_uop_2_stale_dst : _GEN_1345; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1347 = 6'h3 == commit_ptr[5:0] ? rob_uop_3_stale_dst : _GEN_1346; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1348 = 6'h4 == commit_ptr[5:0] ? rob_uop_4_stale_dst : _GEN_1347; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1349 = 6'h5 == commit_ptr[5:0] ? rob_uop_5_stale_dst : _GEN_1348; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1350 = 6'h6 == commit_ptr[5:0] ? rob_uop_6_stale_dst : _GEN_1349; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1351 = 6'h7 == commit_ptr[5:0] ? rob_uop_7_stale_dst : _GEN_1350; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1352 = 6'h8 == commit_ptr[5:0] ? rob_uop_8_stale_dst : _GEN_1351; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1353 = 6'h9 == commit_ptr[5:0] ? rob_uop_9_stale_dst : _GEN_1352; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1354 = 6'ha == commit_ptr[5:0] ? rob_uop_10_stale_dst : _GEN_1353; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1355 = 6'hb == commit_ptr[5:0] ? rob_uop_11_stale_dst : _GEN_1354; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1356 = 6'hc == commit_ptr[5:0] ? rob_uop_12_stale_dst : _GEN_1355; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1357 = 6'hd == commit_ptr[5:0] ? rob_uop_13_stale_dst : _GEN_1356; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1358 = 6'he == commit_ptr[5:0] ? rob_uop_14_stale_dst : _GEN_1357; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1359 = 6'hf == commit_ptr[5:0] ? rob_uop_15_stale_dst : _GEN_1358; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1360 = 6'h10 == commit_ptr[5:0] ? rob_uop_16_stale_dst : _GEN_1359; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1361 = 6'h11 == commit_ptr[5:0] ? rob_uop_17_stale_dst : _GEN_1360; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1362 = 6'h12 == commit_ptr[5:0] ? rob_uop_18_stale_dst : _GEN_1361; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1363 = 6'h13 == commit_ptr[5:0] ? rob_uop_19_stale_dst : _GEN_1362; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1364 = 6'h14 == commit_ptr[5:0] ? rob_uop_20_stale_dst : _GEN_1363; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1365 = 6'h15 == commit_ptr[5:0] ? rob_uop_21_stale_dst : _GEN_1364; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1366 = 6'h16 == commit_ptr[5:0] ? rob_uop_22_stale_dst : _GEN_1365; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1367 = 6'h17 == commit_ptr[5:0] ? rob_uop_23_stale_dst : _GEN_1366; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1368 = 6'h18 == commit_ptr[5:0] ? rob_uop_24_stale_dst : _GEN_1367; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1369 = 6'h19 == commit_ptr[5:0] ? rob_uop_25_stale_dst : _GEN_1368; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1370 = 6'h1a == commit_ptr[5:0] ? rob_uop_26_stale_dst : _GEN_1369; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1371 = 6'h1b == commit_ptr[5:0] ? rob_uop_27_stale_dst : _GEN_1370; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1372 = 6'h1c == commit_ptr[5:0] ? rob_uop_28_stale_dst : _GEN_1371; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1373 = 6'h1d == commit_ptr[5:0] ? rob_uop_29_stale_dst : _GEN_1372; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1374 = 6'h1e == commit_ptr[5:0] ? rob_uop_30_stale_dst : _GEN_1373; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1375 = 6'h1f == commit_ptr[5:0] ? rob_uop_31_stale_dst : _GEN_1374; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1376 = 6'h20 == commit_ptr[5:0] ? rob_uop_32_stale_dst : _GEN_1375; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1377 = 6'h21 == commit_ptr[5:0] ? rob_uop_33_stale_dst : _GEN_1376; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1378 = 6'h22 == commit_ptr[5:0] ? rob_uop_34_stale_dst : _GEN_1377; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1379 = 6'h23 == commit_ptr[5:0] ? rob_uop_35_stale_dst : _GEN_1378; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1380 = 6'h24 == commit_ptr[5:0] ? rob_uop_36_stale_dst : _GEN_1379; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1381 = 6'h25 == commit_ptr[5:0] ? rob_uop_37_stale_dst : _GEN_1380; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1382 = 6'h26 == commit_ptr[5:0] ? rob_uop_38_stale_dst : _GEN_1381; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1383 = 6'h27 == commit_ptr[5:0] ? rob_uop_39_stale_dst : _GEN_1382; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1384 = 6'h28 == commit_ptr[5:0] ? rob_uop_40_stale_dst : _GEN_1383; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1385 = 6'h29 == commit_ptr[5:0] ? rob_uop_41_stale_dst : _GEN_1384; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1386 = 6'h2a == commit_ptr[5:0] ? rob_uop_42_stale_dst : _GEN_1385; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1387 = 6'h2b == commit_ptr[5:0] ? rob_uop_43_stale_dst : _GEN_1386; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1388 = 6'h2c == commit_ptr[5:0] ? rob_uop_44_stale_dst : _GEN_1387; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1389 = 6'h2d == commit_ptr[5:0] ? rob_uop_45_stale_dst : _GEN_1388; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1390 = 6'h2e == commit_ptr[5:0] ? rob_uop_46_stale_dst : _GEN_1389; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1391 = 6'h2f == commit_ptr[5:0] ? rob_uop_47_stale_dst : _GEN_1390; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1392 = 6'h30 == commit_ptr[5:0] ? rob_uop_48_stale_dst : _GEN_1391; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1393 = 6'h31 == commit_ptr[5:0] ? rob_uop_49_stale_dst : _GEN_1392; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1394 = 6'h32 == commit_ptr[5:0] ? rob_uop_50_stale_dst : _GEN_1393; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1395 = 6'h33 == commit_ptr[5:0] ? rob_uop_51_stale_dst : _GEN_1394; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1396 = 6'h34 == commit_ptr[5:0] ? rob_uop_52_stale_dst : _GEN_1395; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1397 = 6'h35 == commit_ptr[5:0] ? rob_uop_53_stale_dst : _GEN_1396; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1398 = 6'h36 == commit_ptr[5:0] ? rob_uop_54_stale_dst : _GEN_1397; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1399 = 6'h37 == commit_ptr[5:0] ? rob_uop_55_stale_dst : _GEN_1398; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1400 = 6'h38 == commit_ptr[5:0] ? rob_uop_56_stale_dst : _GEN_1399; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1401 = 6'h39 == commit_ptr[5:0] ? rob_uop_57_stale_dst : _GEN_1400; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1402 = 6'h3a == commit_ptr[5:0] ? rob_uop_58_stale_dst : _GEN_1401; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1403 = 6'h3b == commit_ptr[5:0] ? rob_uop_59_stale_dst : _GEN_1402; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1404 = 6'h3c == commit_ptr[5:0] ? rob_uop_60_stale_dst : _GEN_1403; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1405 = 6'h3d == commit_ptr[5:0] ? rob_uop_61_stale_dst : _GEN_1404; // @[rob.scala 108:{32,32}]
  wire [6:0] _GEN_1406 = 6'h3e == commit_ptr[5:0] ? rob_uop_62_stale_dst : _GEN_1405; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1409 = 6'h1 == commit_ptr[5:0] ? rob_uop_1_arch_dst : rob_uop_0_arch_dst; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1410 = 6'h2 == commit_ptr[5:0] ? rob_uop_2_arch_dst : _GEN_1409; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1411 = 6'h3 == commit_ptr[5:0] ? rob_uop_3_arch_dst : _GEN_1410; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1412 = 6'h4 == commit_ptr[5:0] ? rob_uop_4_arch_dst : _GEN_1411; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1413 = 6'h5 == commit_ptr[5:0] ? rob_uop_5_arch_dst : _GEN_1412; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1414 = 6'h6 == commit_ptr[5:0] ? rob_uop_6_arch_dst : _GEN_1413; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1415 = 6'h7 == commit_ptr[5:0] ? rob_uop_7_arch_dst : _GEN_1414; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1416 = 6'h8 == commit_ptr[5:0] ? rob_uop_8_arch_dst : _GEN_1415; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1417 = 6'h9 == commit_ptr[5:0] ? rob_uop_9_arch_dst : _GEN_1416; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1418 = 6'ha == commit_ptr[5:0] ? rob_uop_10_arch_dst : _GEN_1417; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1419 = 6'hb == commit_ptr[5:0] ? rob_uop_11_arch_dst : _GEN_1418; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1420 = 6'hc == commit_ptr[5:0] ? rob_uop_12_arch_dst : _GEN_1419; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1421 = 6'hd == commit_ptr[5:0] ? rob_uop_13_arch_dst : _GEN_1420; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1422 = 6'he == commit_ptr[5:0] ? rob_uop_14_arch_dst : _GEN_1421; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1423 = 6'hf == commit_ptr[5:0] ? rob_uop_15_arch_dst : _GEN_1422; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1424 = 6'h10 == commit_ptr[5:0] ? rob_uop_16_arch_dst : _GEN_1423; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1425 = 6'h11 == commit_ptr[5:0] ? rob_uop_17_arch_dst : _GEN_1424; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1426 = 6'h12 == commit_ptr[5:0] ? rob_uop_18_arch_dst : _GEN_1425; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1427 = 6'h13 == commit_ptr[5:0] ? rob_uop_19_arch_dst : _GEN_1426; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1428 = 6'h14 == commit_ptr[5:0] ? rob_uop_20_arch_dst : _GEN_1427; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1429 = 6'h15 == commit_ptr[5:0] ? rob_uop_21_arch_dst : _GEN_1428; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1430 = 6'h16 == commit_ptr[5:0] ? rob_uop_22_arch_dst : _GEN_1429; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1431 = 6'h17 == commit_ptr[5:0] ? rob_uop_23_arch_dst : _GEN_1430; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1432 = 6'h18 == commit_ptr[5:0] ? rob_uop_24_arch_dst : _GEN_1431; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1433 = 6'h19 == commit_ptr[5:0] ? rob_uop_25_arch_dst : _GEN_1432; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1434 = 6'h1a == commit_ptr[5:0] ? rob_uop_26_arch_dst : _GEN_1433; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1435 = 6'h1b == commit_ptr[5:0] ? rob_uop_27_arch_dst : _GEN_1434; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1436 = 6'h1c == commit_ptr[5:0] ? rob_uop_28_arch_dst : _GEN_1435; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1437 = 6'h1d == commit_ptr[5:0] ? rob_uop_29_arch_dst : _GEN_1436; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1438 = 6'h1e == commit_ptr[5:0] ? rob_uop_30_arch_dst : _GEN_1437; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1439 = 6'h1f == commit_ptr[5:0] ? rob_uop_31_arch_dst : _GEN_1438; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1440 = 6'h20 == commit_ptr[5:0] ? rob_uop_32_arch_dst : _GEN_1439; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1441 = 6'h21 == commit_ptr[5:0] ? rob_uop_33_arch_dst : _GEN_1440; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1442 = 6'h22 == commit_ptr[5:0] ? rob_uop_34_arch_dst : _GEN_1441; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1443 = 6'h23 == commit_ptr[5:0] ? rob_uop_35_arch_dst : _GEN_1442; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1444 = 6'h24 == commit_ptr[5:0] ? rob_uop_36_arch_dst : _GEN_1443; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1445 = 6'h25 == commit_ptr[5:0] ? rob_uop_37_arch_dst : _GEN_1444; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1446 = 6'h26 == commit_ptr[5:0] ? rob_uop_38_arch_dst : _GEN_1445; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1447 = 6'h27 == commit_ptr[5:0] ? rob_uop_39_arch_dst : _GEN_1446; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1448 = 6'h28 == commit_ptr[5:0] ? rob_uop_40_arch_dst : _GEN_1447; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1449 = 6'h29 == commit_ptr[5:0] ? rob_uop_41_arch_dst : _GEN_1448; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1450 = 6'h2a == commit_ptr[5:0] ? rob_uop_42_arch_dst : _GEN_1449; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1451 = 6'h2b == commit_ptr[5:0] ? rob_uop_43_arch_dst : _GEN_1450; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1452 = 6'h2c == commit_ptr[5:0] ? rob_uop_44_arch_dst : _GEN_1451; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1453 = 6'h2d == commit_ptr[5:0] ? rob_uop_45_arch_dst : _GEN_1452; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1454 = 6'h2e == commit_ptr[5:0] ? rob_uop_46_arch_dst : _GEN_1453; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1455 = 6'h2f == commit_ptr[5:0] ? rob_uop_47_arch_dst : _GEN_1454; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1456 = 6'h30 == commit_ptr[5:0] ? rob_uop_48_arch_dst : _GEN_1455; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1457 = 6'h31 == commit_ptr[5:0] ? rob_uop_49_arch_dst : _GEN_1456; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1458 = 6'h32 == commit_ptr[5:0] ? rob_uop_50_arch_dst : _GEN_1457; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1459 = 6'h33 == commit_ptr[5:0] ? rob_uop_51_arch_dst : _GEN_1458; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1460 = 6'h34 == commit_ptr[5:0] ? rob_uop_52_arch_dst : _GEN_1459; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1461 = 6'h35 == commit_ptr[5:0] ? rob_uop_53_arch_dst : _GEN_1460; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1462 = 6'h36 == commit_ptr[5:0] ? rob_uop_54_arch_dst : _GEN_1461; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1463 = 6'h37 == commit_ptr[5:0] ? rob_uop_55_arch_dst : _GEN_1462; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1464 = 6'h38 == commit_ptr[5:0] ? rob_uop_56_arch_dst : _GEN_1463; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1465 = 6'h39 == commit_ptr[5:0] ? rob_uop_57_arch_dst : _GEN_1464; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1466 = 6'h3a == commit_ptr[5:0] ? rob_uop_58_arch_dst : _GEN_1465; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1467 = 6'h3b == commit_ptr[5:0] ? rob_uop_59_arch_dst : _GEN_1466; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1468 = 6'h3c == commit_ptr[5:0] ? rob_uop_60_arch_dst : _GEN_1467; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1469 = 6'h3d == commit_ptr[5:0] ? rob_uop_61_arch_dst : _GEN_1468; // @[rob.scala 108:{32,32}]
  wire [4:0] _GEN_1470 = 6'h3e == commit_ptr[5:0] ? rob_uop_62_arch_dst : _GEN_1469; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2113 = 6'h1 == commit_ptr[5:0] ? rob_uop_1_dst_value : rob_uop_0_dst_value; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2114 = 6'h2 == commit_ptr[5:0] ? rob_uop_2_dst_value : _GEN_2113; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2115 = 6'h3 == commit_ptr[5:0] ? rob_uop_3_dst_value : _GEN_2114; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2116 = 6'h4 == commit_ptr[5:0] ? rob_uop_4_dst_value : _GEN_2115; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2117 = 6'h5 == commit_ptr[5:0] ? rob_uop_5_dst_value : _GEN_2116; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2118 = 6'h6 == commit_ptr[5:0] ? rob_uop_6_dst_value : _GEN_2117; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2119 = 6'h7 == commit_ptr[5:0] ? rob_uop_7_dst_value : _GEN_2118; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2120 = 6'h8 == commit_ptr[5:0] ? rob_uop_8_dst_value : _GEN_2119; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2121 = 6'h9 == commit_ptr[5:0] ? rob_uop_9_dst_value : _GEN_2120; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2122 = 6'ha == commit_ptr[5:0] ? rob_uop_10_dst_value : _GEN_2121; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2123 = 6'hb == commit_ptr[5:0] ? rob_uop_11_dst_value : _GEN_2122; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2124 = 6'hc == commit_ptr[5:0] ? rob_uop_12_dst_value : _GEN_2123; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2125 = 6'hd == commit_ptr[5:0] ? rob_uop_13_dst_value : _GEN_2124; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2126 = 6'he == commit_ptr[5:0] ? rob_uop_14_dst_value : _GEN_2125; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2127 = 6'hf == commit_ptr[5:0] ? rob_uop_15_dst_value : _GEN_2126; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2128 = 6'h10 == commit_ptr[5:0] ? rob_uop_16_dst_value : _GEN_2127; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2129 = 6'h11 == commit_ptr[5:0] ? rob_uop_17_dst_value : _GEN_2128; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2130 = 6'h12 == commit_ptr[5:0] ? rob_uop_18_dst_value : _GEN_2129; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2131 = 6'h13 == commit_ptr[5:0] ? rob_uop_19_dst_value : _GEN_2130; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2132 = 6'h14 == commit_ptr[5:0] ? rob_uop_20_dst_value : _GEN_2131; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2133 = 6'h15 == commit_ptr[5:0] ? rob_uop_21_dst_value : _GEN_2132; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2134 = 6'h16 == commit_ptr[5:0] ? rob_uop_22_dst_value : _GEN_2133; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2135 = 6'h17 == commit_ptr[5:0] ? rob_uop_23_dst_value : _GEN_2134; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2136 = 6'h18 == commit_ptr[5:0] ? rob_uop_24_dst_value : _GEN_2135; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2137 = 6'h19 == commit_ptr[5:0] ? rob_uop_25_dst_value : _GEN_2136; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2138 = 6'h1a == commit_ptr[5:0] ? rob_uop_26_dst_value : _GEN_2137; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2139 = 6'h1b == commit_ptr[5:0] ? rob_uop_27_dst_value : _GEN_2138; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2140 = 6'h1c == commit_ptr[5:0] ? rob_uop_28_dst_value : _GEN_2139; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2141 = 6'h1d == commit_ptr[5:0] ? rob_uop_29_dst_value : _GEN_2140; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2142 = 6'h1e == commit_ptr[5:0] ? rob_uop_30_dst_value : _GEN_2141; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2143 = 6'h1f == commit_ptr[5:0] ? rob_uop_31_dst_value : _GEN_2142; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2144 = 6'h20 == commit_ptr[5:0] ? rob_uop_32_dst_value : _GEN_2143; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2145 = 6'h21 == commit_ptr[5:0] ? rob_uop_33_dst_value : _GEN_2144; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2146 = 6'h22 == commit_ptr[5:0] ? rob_uop_34_dst_value : _GEN_2145; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2147 = 6'h23 == commit_ptr[5:0] ? rob_uop_35_dst_value : _GEN_2146; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2148 = 6'h24 == commit_ptr[5:0] ? rob_uop_36_dst_value : _GEN_2147; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2149 = 6'h25 == commit_ptr[5:0] ? rob_uop_37_dst_value : _GEN_2148; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2150 = 6'h26 == commit_ptr[5:0] ? rob_uop_38_dst_value : _GEN_2149; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2151 = 6'h27 == commit_ptr[5:0] ? rob_uop_39_dst_value : _GEN_2150; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2152 = 6'h28 == commit_ptr[5:0] ? rob_uop_40_dst_value : _GEN_2151; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2153 = 6'h29 == commit_ptr[5:0] ? rob_uop_41_dst_value : _GEN_2152; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2154 = 6'h2a == commit_ptr[5:0] ? rob_uop_42_dst_value : _GEN_2153; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2155 = 6'h2b == commit_ptr[5:0] ? rob_uop_43_dst_value : _GEN_2154; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2156 = 6'h2c == commit_ptr[5:0] ? rob_uop_44_dst_value : _GEN_2155; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2157 = 6'h2d == commit_ptr[5:0] ? rob_uop_45_dst_value : _GEN_2156; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2158 = 6'h2e == commit_ptr[5:0] ? rob_uop_46_dst_value : _GEN_2157; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2159 = 6'h2f == commit_ptr[5:0] ? rob_uop_47_dst_value : _GEN_2158; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2160 = 6'h30 == commit_ptr[5:0] ? rob_uop_48_dst_value : _GEN_2159; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2161 = 6'h31 == commit_ptr[5:0] ? rob_uop_49_dst_value : _GEN_2160; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2162 = 6'h32 == commit_ptr[5:0] ? rob_uop_50_dst_value : _GEN_2161; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2163 = 6'h33 == commit_ptr[5:0] ? rob_uop_51_dst_value : _GEN_2162; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2164 = 6'h34 == commit_ptr[5:0] ? rob_uop_52_dst_value : _GEN_2163; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2165 = 6'h35 == commit_ptr[5:0] ? rob_uop_53_dst_value : _GEN_2164; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2166 = 6'h36 == commit_ptr[5:0] ? rob_uop_54_dst_value : _GEN_2165; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2167 = 6'h37 == commit_ptr[5:0] ? rob_uop_55_dst_value : _GEN_2166; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2168 = 6'h38 == commit_ptr[5:0] ? rob_uop_56_dst_value : _GEN_2167; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2169 = 6'h39 == commit_ptr[5:0] ? rob_uop_57_dst_value : _GEN_2168; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2170 = 6'h3a == commit_ptr[5:0] ? rob_uop_58_dst_value : _GEN_2169; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2171 = 6'h3b == commit_ptr[5:0] ? rob_uop_59_dst_value : _GEN_2170; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2172 = 6'h3c == commit_ptr[5:0] ? rob_uop_60_dst_value : _GEN_2171; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2173 = 6'h3d == commit_ptr[5:0] ? rob_uop_61_dst_value : _GEN_2172; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2174 = 6'h3e == commit_ptr[5:0] ? rob_uop_62_dst_value : _GEN_2173; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2177 = 6'h1 == commit_ptr[5:0] ? rob_uop_1_src1_value : rob_uop_0_src1_value; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2178 = 6'h2 == commit_ptr[5:0] ? rob_uop_2_src1_value : _GEN_2177; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2179 = 6'h3 == commit_ptr[5:0] ? rob_uop_3_src1_value : _GEN_2178; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2180 = 6'h4 == commit_ptr[5:0] ? rob_uop_4_src1_value : _GEN_2179; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2181 = 6'h5 == commit_ptr[5:0] ? rob_uop_5_src1_value : _GEN_2180; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2182 = 6'h6 == commit_ptr[5:0] ? rob_uop_6_src1_value : _GEN_2181; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2183 = 6'h7 == commit_ptr[5:0] ? rob_uop_7_src1_value : _GEN_2182; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2184 = 6'h8 == commit_ptr[5:0] ? rob_uop_8_src1_value : _GEN_2183; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2185 = 6'h9 == commit_ptr[5:0] ? rob_uop_9_src1_value : _GEN_2184; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2186 = 6'ha == commit_ptr[5:0] ? rob_uop_10_src1_value : _GEN_2185; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2187 = 6'hb == commit_ptr[5:0] ? rob_uop_11_src1_value : _GEN_2186; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2188 = 6'hc == commit_ptr[5:0] ? rob_uop_12_src1_value : _GEN_2187; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2189 = 6'hd == commit_ptr[5:0] ? rob_uop_13_src1_value : _GEN_2188; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2190 = 6'he == commit_ptr[5:0] ? rob_uop_14_src1_value : _GEN_2189; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2191 = 6'hf == commit_ptr[5:0] ? rob_uop_15_src1_value : _GEN_2190; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2192 = 6'h10 == commit_ptr[5:0] ? rob_uop_16_src1_value : _GEN_2191; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2193 = 6'h11 == commit_ptr[5:0] ? rob_uop_17_src1_value : _GEN_2192; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2194 = 6'h12 == commit_ptr[5:0] ? rob_uop_18_src1_value : _GEN_2193; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2195 = 6'h13 == commit_ptr[5:0] ? rob_uop_19_src1_value : _GEN_2194; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2196 = 6'h14 == commit_ptr[5:0] ? rob_uop_20_src1_value : _GEN_2195; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2197 = 6'h15 == commit_ptr[5:0] ? rob_uop_21_src1_value : _GEN_2196; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2198 = 6'h16 == commit_ptr[5:0] ? rob_uop_22_src1_value : _GEN_2197; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2199 = 6'h17 == commit_ptr[5:0] ? rob_uop_23_src1_value : _GEN_2198; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2200 = 6'h18 == commit_ptr[5:0] ? rob_uop_24_src1_value : _GEN_2199; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2201 = 6'h19 == commit_ptr[5:0] ? rob_uop_25_src1_value : _GEN_2200; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2202 = 6'h1a == commit_ptr[5:0] ? rob_uop_26_src1_value : _GEN_2201; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2203 = 6'h1b == commit_ptr[5:0] ? rob_uop_27_src1_value : _GEN_2202; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2204 = 6'h1c == commit_ptr[5:0] ? rob_uop_28_src1_value : _GEN_2203; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2205 = 6'h1d == commit_ptr[5:0] ? rob_uop_29_src1_value : _GEN_2204; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2206 = 6'h1e == commit_ptr[5:0] ? rob_uop_30_src1_value : _GEN_2205; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2207 = 6'h1f == commit_ptr[5:0] ? rob_uop_31_src1_value : _GEN_2206; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2208 = 6'h20 == commit_ptr[5:0] ? rob_uop_32_src1_value : _GEN_2207; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2209 = 6'h21 == commit_ptr[5:0] ? rob_uop_33_src1_value : _GEN_2208; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2210 = 6'h22 == commit_ptr[5:0] ? rob_uop_34_src1_value : _GEN_2209; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2211 = 6'h23 == commit_ptr[5:0] ? rob_uop_35_src1_value : _GEN_2210; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2212 = 6'h24 == commit_ptr[5:0] ? rob_uop_36_src1_value : _GEN_2211; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2213 = 6'h25 == commit_ptr[5:0] ? rob_uop_37_src1_value : _GEN_2212; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2214 = 6'h26 == commit_ptr[5:0] ? rob_uop_38_src1_value : _GEN_2213; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2215 = 6'h27 == commit_ptr[5:0] ? rob_uop_39_src1_value : _GEN_2214; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2216 = 6'h28 == commit_ptr[5:0] ? rob_uop_40_src1_value : _GEN_2215; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2217 = 6'h29 == commit_ptr[5:0] ? rob_uop_41_src1_value : _GEN_2216; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2218 = 6'h2a == commit_ptr[5:0] ? rob_uop_42_src1_value : _GEN_2217; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2219 = 6'h2b == commit_ptr[5:0] ? rob_uop_43_src1_value : _GEN_2218; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2220 = 6'h2c == commit_ptr[5:0] ? rob_uop_44_src1_value : _GEN_2219; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2221 = 6'h2d == commit_ptr[5:0] ? rob_uop_45_src1_value : _GEN_2220; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2222 = 6'h2e == commit_ptr[5:0] ? rob_uop_46_src1_value : _GEN_2221; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2223 = 6'h2f == commit_ptr[5:0] ? rob_uop_47_src1_value : _GEN_2222; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2224 = 6'h30 == commit_ptr[5:0] ? rob_uop_48_src1_value : _GEN_2223; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2225 = 6'h31 == commit_ptr[5:0] ? rob_uop_49_src1_value : _GEN_2224; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2226 = 6'h32 == commit_ptr[5:0] ? rob_uop_50_src1_value : _GEN_2225; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2227 = 6'h33 == commit_ptr[5:0] ? rob_uop_51_src1_value : _GEN_2226; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2228 = 6'h34 == commit_ptr[5:0] ? rob_uop_52_src1_value : _GEN_2227; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2229 = 6'h35 == commit_ptr[5:0] ? rob_uop_53_src1_value : _GEN_2228; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2230 = 6'h36 == commit_ptr[5:0] ? rob_uop_54_src1_value : _GEN_2229; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2231 = 6'h37 == commit_ptr[5:0] ? rob_uop_55_src1_value : _GEN_2230; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2232 = 6'h38 == commit_ptr[5:0] ? rob_uop_56_src1_value : _GEN_2231; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2233 = 6'h39 == commit_ptr[5:0] ? rob_uop_57_src1_value : _GEN_2232; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2234 = 6'h3a == commit_ptr[5:0] ? rob_uop_58_src1_value : _GEN_2233; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2235 = 6'h3b == commit_ptr[5:0] ? rob_uop_59_src1_value : _GEN_2234; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2236 = 6'h3c == commit_ptr[5:0] ? rob_uop_60_src1_value : _GEN_2235; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2237 = 6'h3d == commit_ptr[5:0] ? rob_uop_61_src1_value : _GEN_2236; // @[rob.scala 108:{32,32}]
  wire [63:0] _GEN_2238 = 6'h3e == commit_ptr[5:0] ? rob_uop_62_src1_value : _GEN_2237; // @[rob.scala 108:{32,32}]
  wire [31:0] _GEN_2817 = 6'h1 == _next_can_commit_1_T_1[5:0] ? rob_uop_1_inst : rob_uop_0_inst; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2818 = 6'h2 == _next_can_commit_1_T_1[5:0] ? rob_uop_2_inst : _GEN_2817; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2819 = 6'h3 == _next_can_commit_1_T_1[5:0] ? rob_uop_3_inst : _GEN_2818; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2820 = 6'h4 == _next_can_commit_1_T_1[5:0] ? rob_uop_4_inst : _GEN_2819; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2821 = 6'h5 == _next_can_commit_1_T_1[5:0] ? rob_uop_5_inst : _GEN_2820; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2822 = 6'h6 == _next_can_commit_1_T_1[5:0] ? rob_uop_6_inst : _GEN_2821; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2823 = 6'h7 == _next_can_commit_1_T_1[5:0] ? rob_uop_7_inst : _GEN_2822; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2824 = 6'h8 == _next_can_commit_1_T_1[5:0] ? rob_uop_8_inst : _GEN_2823; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2825 = 6'h9 == _next_can_commit_1_T_1[5:0] ? rob_uop_9_inst : _GEN_2824; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2826 = 6'ha == _next_can_commit_1_T_1[5:0] ? rob_uop_10_inst : _GEN_2825; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2827 = 6'hb == _next_can_commit_1_T_1[5:0] ? rob_uop_11_inst : _GEN_2826; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2828 = 6'hc == _next_can_commit_1_T_1[5:0] ? rob_uop_12_inst : _GEN_2827; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2829 = 6'hd == _next_can_commit_1_T_1[5:0] ? rob_uop_13_inst : _GEN_2828; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2830 = 6'he == _next_can_commit_1_T_1[5:0] ? rob_uop_14_inst : _GEN_2829; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2831 = 6'hf == _next_can_commit_1_T_1[5:0] ? rob_uop_15_inst : _GEN_2830; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2832 = 6'h10 == _next_can_commit_1_T_1[5:0] ? rob_uop_16_inst : _GEN_2831; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2833 = 6'h11 == _next_can_commit_1_T_1[5:0] ? rob_uop_17_inst : _GEN_2832; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2834 = 6'h12 == _next_can_commit_1_T_1[5:0] ? rob_uop_18_inst : _GEN_2833; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2835 = 6'h13 == _next_can_commit_1_T_1[5:0] ? rob_uop_19_inst : _GEN_2834; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2836 = 6'h14 == _next_can_commit_1_T_1[5:0] ? rob_uop_20_inst : _GEN_2835; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2837 = 6'h15 == _next_can_commit_1_T_1[5:0] ? rob_uop_21_inst : _GEN_2836; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2838 = 6'h16 == _next_can_commit_1_T_1[5:0] ? rob_uop_22_inst : _GEN_2837; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2839 = 6'h17 == _next_can_commit_1_T_1[5:0] ? rob_uop_23_inst : _GEN_2838; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2840 = 6'h18 == _next_can_commit_1_T_1[5:0] ? rob_uop_24_inst : _GEN_2839; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2841 = 6'h19 == _next_can_commit_1_T_1[5:0] ? rob_uop_25_inst : _GEN_2840; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2842 = 6'h1a == _next_can_commit_1_T_1[5:0] ? rob_uop_26_inst : _GEN_2841; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2843 = 6'h1b == _next_can_commit_1_T_1[5:0] ? rob_uop_27_inst : _GEN_2842; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2844 = 6'h1c == _next_can_commit_1_T_1[5:0] ? rob_uop_28_inst : _GEN_2843; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2845 = 6'h1d == _next_can_commit_1_T_1[5:0] ? rob_uop_29_inst : _GEN_2844; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2846 = 6'h1e == _next_can_commit_1_T_1[5:0] ? rob_uop_30_inst : _GEN_2845; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2847 = 6'h1f == _next_can_commit_1_T_1[5:0] ? rob_uop_31_inst : _GEN_2846; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2848 = 6'h20 == _next_can_commit_1_T_1[5:0] ? rob_uop_32_inst : _GEN_2847; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2849 = 6'h21 == _next_can_commit_1_T_1[5:0] ? rob_uop_33_inst : _GEN_2848; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2850 = 6'h22 == _next_can_commit_1_T_1[5:0] ? rob_uop_34_inst : _GEN_2849; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2851 = 6'h23 == _next_can_commit_1_T_1[5:0] ? rob_uop_35_inst : _GEN_2850; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2852 = 6'h24 == _next_can_commit_1_T_1[5:0] ? rob_uop_36_inst : _GEN_2851; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2853 = 6'h25 == _next_can_commit_1_T_1[5:0] ? rob_uop_37_inst : _GEN_2852; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2854 = 6'h26 == _next_can_commit_1_T_1[5:0] ? rob_uop_38_inst : _GEN_2853; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2855 = 6'h27 == _next_can_commit_1_T_1[5:0] ? rob_uop_39_inst : _GEN_2854; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2856 = 6'h28 == _next_can_commit_1_T_1[5:0] ? rob_uop_40_inst : _GEN_2855; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2857 = 6'h29 == _next_can_commit_1_T_1[5:0] ? rob_uop_41_inst : _GEN_2856; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2858 = 6'h2a == _next_can_commit_1_T_1[5:0] ? rob_uop_42_inst : _GEN_2857; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2859 = 6'h2b == _next_can_commit_1_T_1[5:0] ? rob_uop_43_inst : _GEN_2858; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2860 = 6'h2c == _next_can_commit_1_T_1[5:0] ? rob_uop_44_inst : _GEN_2859; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2861 = 6'h2d == _next_can_commit_1_T_1[5:0] ? rob_uop_45_inst : _GEN_2860; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2862 = 6'h2e == _next_can_commit_1_T_1[5:0] ? rob_uop_46_inst : _GEN_2861; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2863 = 6'h2f == _next_can_commit_1_T_1[5:0] ? rob_uop_47_inst : _GEN_2862; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2864 = 6'h30 == _next_can_commit_1_T_1[5:0] ? rob_uop_48_inst : _GEN_2863; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2865 = 6'h31 == _next_can_commit_1_T_1[5:0] ? rob_uop_49_inst : _GEN_2864; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2866 = 6'h32 == _next_can_commit_1_T_1[5:0] ? rob_uop_50_inst : _GEN_2865; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2867 = 6'h33 == _next_can_commit_1_T_1[5:0] ? rob_uop_51_inst : _GEN_2866; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2868 = 6'h34 == _next_can_commit_1_T_1[5:0] ? rob_uop_52_inst : _GEN_2867; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2869 = 6'h35 == _next_can_commit_1_T_1[5:0] ? rob_uop_53_inst : _GEN_2868; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2870 = 6'h36 == _next_can_commit_1_T_1[5:0] ? rob_uop_54_inst : _GEN_2869; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2871 = 6'h37 == _next_can_commit_1_T_1[5:0] ? rob_uop_55_inst : _GEN_2870; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2872 = 6'h38 == _next_can_commit_1_T_1[5:0] ? rob_uop_56_inst : _GEN_2871; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2873 = 6'h39 == _next_can_commit_1_T_1[5:0] ? rob_uop_57_inst : _GEN_2872; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2874 = 6'h3a == _next_can_commit_1_T_1[5:0] ? rob_uop_58_inst : _GEN_2873; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2875 = 6'h3b == _next_can_commit_1_T_1[5:0] ? rob_uop_59_inst : _GEN_2874; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2876 = 6'h3c == _next_can_commit_1_T_1[5:0] ? rob_uop_60_inst : _GEN_2875; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2877 = 6'h3d == _next_can_commit_1_T_1[5:0] ? rob_uop_61_inst : _GEN_2876; // @[rob.scala 109:{32,32}]
  wire [31:0] _GEN_2878 = 6'h3e == _next_can_commit_1_T_1[5:0] ? rob_uop_62_inst : _GEN_2877; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2881 = 6'h1 == _next_can_commit_1_T_1[5:0] ? rob_uop_1_func_code : rob_uop_0_func_code; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2882 = 6'h2 == _next_can_commit_1_T_1[5:0] ? rob_uop_2_func_code : _GEN_2881; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2883 = 6'h3 == _next_can_commit_1_T_1[5:0] ? rob_uop_3_func_code : _GEN_2882; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2884 = 6'h4 == _next_can_commit_1_T_1[5:0] ? rob_uop_4_func_code : _GEN_2883; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2885 = 6'h5 == _next_can_commit_1_T_1[5:0] ? rob_uop_5_func_code : _GEN_2884; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2886 = 6'h6 == _next_can_commit_1_T_1[5:0] ? rob_uop_6_func_code : _GEN_2885; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2887 = 6'h7 == _next_can_commit_1_T_1[5:0] ? rob_uop_7_func_code : _GEN_2886; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2888 = 6'h8 == _next_can_commit_1_T_1[5:0] ? rob_uop_8_func_code : _GEN_2887; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2889 = 6'h9 == _next_can_commit_1_T_1[5:0] ? rob_uop_9_func_code : _GEN_2888; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2890 = 6'ha == _next_can_commit_1_T_1[5:0] ? rob_uop_10_func_code : _GEN_2889; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2891 = 6'hb == _next_can_commit_1_T_1[5:0] ? rob_uop_11_func_code : _GEN_2890; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2892 = 6'hc == _next_can_commit_1_T_1[5:0] ? rob_uop_12_func_code : _GEN_2891; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2893 = 6'hd == _next_can_commit_1_T_1[5:0] ? rob_uop_13_func_code : _GEN_2892; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2894 = 6'he == _next_can_commit_1_T_1[5:0] ? rob_uop_14_func_code : _GEN_2893; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2895 = 6'hf == _next_can_commit_1_T_1[5:0] ? rob_uop_15_func_code : _GEN_2894; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2896 = 6'h10 == _next_can_commit_1_T_1[5:0] ? rob_uop_16_func_code : _GEN_2895; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2897 = 6'h11 == _next_can_commit_1_T_1[5:0] ? rob_uop_17_func_code : _GEN_2896; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2898 = 6'h12 == _next_can_commit_1_T_1[5:0] ? rob_uop_18_func_code : _GEN_2897; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2899 = 6'h13 == _next_can_commit_1_T_1[5:0] ? rob_uop_19_func_code : _GEN_2898; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2900 = 6'h14 == _next_can_commit_1_T_1[5:0] ? rob_uop_20_func_code : _GEN_2899; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2901 = 6'h15 == _next_can_commit_1_T_1[5:0] ? rob_uop_21_func_code : _GEN_2900; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2902 = 6'h16 == _next_can_commit_1_T_1[5:0] ? rob_uop_22_func_code : _GEN_2901; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2903 = 6'h17 == _next_can_commit_1_T_1[5:0] ? rob_uop_23_func_code : _GEN_2902; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2904 = 6'h18 == _next_can_commit_1_T_1[5:0] ? rob_uop_24_func_code : _GEN_2903; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2905 = 6'h19 == _next_can_commit_1_T_1[5:0] ? rob_uop_25_func_code : _GEN_2904; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2906 = 6'h1a == _next_can_commit_1_T_1[5:0] ? rob_uop_26_func_code : _GEN_2905; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2907 = 6'h1b == _next_can_commit_1_T_1[5:0] ? rob_uop_27_func_code : _GEN_2906; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2908 = 6'h1c == _next_can_commit_1_T_1[5:0] ? rob_uop_28_func_code : _GEN_2907; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2909 = 6'h1d == _next_can_commit_1_T_1[5:0] ? rob_uop_29_func_code : _GEN_2908; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2910 = 6'h1e == _next_can_commit_1_T_1[5:0] ? rob_uop_30_func_code : _GEN_2909; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2911 = 6'h1f == _next_can_commit_1_T_1[5:0] ? rob_uop_31_func_code : _GEN_2910; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2912 = 6'h20 == _next_can_commit_1_T_1[5:0] ? rob_uop_32_func_code : _GEN_2911; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2913 = 6'h21 == _next_can_commit_1_T_1[5:0] ? rob_uop_33_func_code : _GEN_2912; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2914 = 6'h22 == _next_can_commit_1_T_1[5:0] ? rob_uop_34_func_code : _GEN_2913; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2915 = 6'h23 == _next_can_commit_1_T_1[5:0] ? rob_uop_35_func_code : _GEN_2914; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2916 = 6'h24 == _next_can_commit_1_T_1[5:0] ? rob_uop_36_func_code : _GEN_2915; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2917 = 6'h25 == _next_can_commit_1_T_1[5:0] ? rob_uop_37_func_code : _GEN_2916; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2918 = 6'h26 == _next_can_commit_1_T_1[5:0] ? rob_uop_38_func_code : _GEN_2917; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2919 = 6'h27 == _next_can_commit_1_T_1[5:0] ? rob_uop_39_func_code : _GEN_2918; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2920 = 6'h28 == _next_can_commit_1_T_1[5:0] ? rob_uop_40_func_code : _GEN_2919; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2921 = 6'h29 == _next_can_commit_1_T_1[5:0] ? rob_uop_41_func_code : _GEN_2920; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2922 = 6'h2a == _next_can_commit_1_T_1[5:0] ? rob_uop_42_func_code : _GEN_2921; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2923 = 6'h2b == _next_can_commit_1_T_1[5:0] ? rob_uop_43_func_code : _GEN_2922; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2924 = 6'h2c == _next_can_commit_1_T_1[5:0] ? rob_uop_44_func_code : _GEN_2923; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2925 = 6'h2d == _next_can_commit_1_T_1[5:0] ? rob_uop_45_func_code : _GEN_2924; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2926 = 6'h2e == _next_can_commit_1_T_1[5:0] ? rob_uop_46_func_code : _GEN_2925; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2927 = 6'h2f == _next_can_commit_1_T_1[5:0] ? rob_uop_47_func_code : _GEN_2926; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2928 = 6'h30 == _next_can_commit_1_T_1[5:0] ? rob_uop_48_func_code : _GEN_2927; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2929 = 6'h31 == _next_can_commit_1_T_1[5:0] ? rob_uop_49_func_code : _GEN_2928; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2930 = 6'h32 == _next_can_commit_1_T_1[5:0] ? rob_uop_50_func_code : _GEN_2929; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2931 = 6'h33 == _next_can_commit_1_T_1[5:0] ? rob_uop_51_func_code : _GEN_2930; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2932 = 6'h34 == _next_can_commit_1_T_1[5:0] ? rob_uop_52_func_code : _GEN_2931; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2933 = 6'h35 == _next_can_commit_1_T_1[5:0] ? rob_uop_53_func_code : _GEN_2932; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2934 = 6'h36 == _next_can_commit_1_T_1[5:0] ? rob_uop_54_func_code : _GEN_2933; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2935 = 6'h37 == _next_can_commit_1_T_1[5:0] ? rob_uop_55_func_code : _GEN_2934; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2936 = 6'h38 == _next_can_commit_1_T_1[5:0] ? rob_uop_56_func_code : _GEN_2935; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2937 = 6'h39 == _next_can_commit_1_T_1[5:0] ? rob_uop_57_func_code : _GEN_2936; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2938 = 6'h3a == _next_can_commit_1_T_1[5:0] ? rob_uop_58_func_code : _GEN_2937; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2939 = 6'h3b == _next_can_commit_1_T_1[5:0] ? rob_uop_59_func_code : _GEN_2938; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2940 = 6'h3c == _next_can_commit_1_T_1[5:0] ? rob_uop_60_func_code : _GEN_2939; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2941 = 6'h3d == _next_can_commit_1_T_1[5:0] ? rob_uop_61_func_code : _GEN_2940; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_2942 = 6'h3e == _next_can_commit_1_T_1[5:0] ? rob_uop_62_func_code : _GEN_2941; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3265 = 6'h1 == _next_can_commit_1_T_1[5:0] ? rob_uop_1_phy_dst : rob_uop_0_phy_dst; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3266 = 6'h2 == _next_can_commit_1_T_1[5:0] ? rob_uop_2_phy_dst : _GEN_3265; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3267 = 6'h3 == _next_can_commit_1_T_1[5:0] ? rob_uop_3_phy_dst : _GEN_3266; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3268 = 6'h4 == _next_can_commit_1_T_1[5:0] ? rob_uop_4_phy_dst : _GEN_3267; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3269 = 6'h5 == _next_can_commit_1_T_1[5:0] ? rob_uop_5_phy_dst : _GEN_3268; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3270 = 6'h6 == _next_can_commit_1_T_1[5:0] ? rob_uop_6_phy_dst : _GEN_3269; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3271 = 6'h7 == _next_can_commit_1_T_1[5:0] ? rob_uop_7_phy_dst : _GEN_3270; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3272 = 6'h8 == _next_can_commit_1_T_1[5:0] ? rob_uop_8_phy_dst : _GEN_3271; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3273 = 6'h9 == _next_can_commit_1_T_1[5:0] ? rob_uop_9_phy_dst : _GEN_3272; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3274 = 6'ha == _next_can_commit_1_T_1[5:0] ? rob_uop_10_phy_dst : _GEN_3273; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3275 = 6'hb == _next_can_commit_1_T_1[5:0] ? rob_uop_11_phy_dst : _GEN_3274; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3276 = 6'hc == _next_can_commit_1_T_1[5:0] ? rob_uop_12_phy_dst : _GEN_3275; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3277 = 6'hd == _next_can_commit_1_T_1[5:0] ? rob_uop_13_phy_dst : _GEN_3276; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3278 = 6'he == _next_can_commit_1_T_1[5:0] ? rob_uop_14_phy_dst : _GEN_3277; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3279 = 6'hf == _next_can_commit_1_T_1[5:0] ? rob_uop_15_phy_dst : _GEN_3278; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3280 = 6'h10 == _next_can_commit_1_T_1[5:0] ? rob_uop_16_phy_dst : _GEN_3279; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3281 = 6'h11 == _next_can_commit_1_T_1[5:0] ? rob_uop_17_phy_dst : _GEN_3280; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3282 = 6'h12 == _next_can_commit_1_T_1[5:0] ? rob_uop_18_phy_dst : _GEN_3281; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3283 = 6'h13 == _next_can_commit_1_T_1[5:0] ? rob_uop_19_phy_dst : _GEN_3282; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3284 = 6'h14 == _next_can_commit_1_T_1[5:0] ? rob_uop_20_phy_dst : _GEN_3283; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3285 = 6'h15 == _next_can_commit_1_T_1[5:0] ? rob_uop_21_phy_dst : _GEN_3284; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3286 = 6'h16 == _next_can_commit_1_T_1[5:0] ? rob_uop_22_phy_dst : _GEN_3285; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3287 = 6'h17 == _next_can_commit_1_T_1[5:0] ? rob_uop_23_phy_dst : _GEN_3286; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3288 = 6'h18 == _next_can_commit_1_T_1[5:0] ? rob_uop_24_phy_dst : _GEN_3287; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3289 = 6'h19 == _next_can_commit_1_T_1[5:0] ? rob_uop_25_phy_dst : _GEN_3288; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3290 = 6'h1a == _next_can_commit_1_T_1[5:0] ? rob_uop_26_phy_dst : _GEN_3289; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3291 = 6'h1b == _next_can_commit_1_T_1[5:0] ? rob_uop_27_phy_dst : _GEN_3290; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3292 = 6'h1c == _next_can_commit_1_T_1[5:0] ? rob_uop_28_phy_dst : _GEN_3291; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3293 = 6'h1d == _next_can_commit_1_T_1[5:0] ? rob_uop_29_phy_dst : _GEN_3292; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3294 = 6'h1e == _next_can_commit_1_T_1[5:0] ? rob_uop_30_phy_dst : _GEN_3293; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3295 = 6'h1f == _next_can_commit_1_T_1[5:0] ? rob_uop_31_phy_dst : _GEN_3294; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3296 = 6'h20 == _next_can_commit_1_T_1[5:0] ? rob_uop_32_phy_dst : _GEN_3295; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3297 = 6'h21 == _next_can_commit_1_T_1[5:0] ? rob_uop_33_phy_dst : _GEN_3296; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3298 = 6'h22 == _next_can_commit_1_T_1[5:0] ? rob_uop_34_phy_dst : _GEN_3297; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3299 = 6'h23 == _next_can_commit_1_T_1[5:0] ? rob_uop_35_phy_dst : _GEN_3298; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3300 = 6'h24 == _next_can_commit_1_T_1[5:0] ? rob_uop_36_phy_dst : _GEN_3299; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3301 = 6'h25 == _next_can_commit_1_T_1[5:0] ? rob_uop_37_phy_dst : _GEN_3300; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3302 = 6'h26 == _next_can_commit_1_T_1[5:0] ? rob_uop_38_phy_dst : _GEN_3301; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3303 = 6'h27 == _next_can_commit_1_T_1[5:0] ? rob_uop_39_phy_dst : _GEN_3302; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3304 = 6'h28 == _next_can_commit_1_T_1[5:0] ? rob_uop_40_phy_dst : _GEN_3303; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3305 = 6'h29 == _next_can_commit_1_T_1[5:0] ? rob_uop_41_phy_dst : _GEN_3304; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3306 = 6'h2a == _next_can_commit_1_T_1[5:0] ? rob_uop_42_phy_dst : _GEN_3305; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3307 = 6'h2b == _next_can_commit_1_T_1[5:0] ? rob_uop_43_phy_dst : _GEN_3306; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3308 = 6'h2c == _next_can_commit_1_T_1[5:0] ? rob_uop_44_phy_dst : _GEN_3307; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3309 = 6'h2d == _next_can_commit_1_T_1[5:0] ? rob_uop_45_phy_dst : _GEN_3308; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3310 = 6'h2e == _next_can_commit_1_T_1[5:0] ? rob_uop_46_phy_dst : _GEN_3309; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3311 = 6'h2f == _next_can_commit_1_T_1[5:0] ? rob_uop_47_phy_dst : _GEN_3310; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3312 = 6'h30 == _next_can_commit_1_T_1[5:0] ? rob_uop_48_phy_dst : _GEN_3311; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3313 = 6'h31 == _next_can_commit_1_T_1[5:0] ? rob_uop_49_phy_dst : _GEN_3312; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3314 = 6'h32 == _next_can_commit_1_T_1[5:0] ? rob_uop_50_phy_dst : _GEN_3313; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3315 = 6'h33 == _next_can_commit_1_T_1[5:0] ? rob_uop_51_phy_dst : _GEN_3314; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3316 = 6'h34 == _next_can_commit_1_T_1[5:0] ? rob_uop_52_phy_dst : _GEN_3315; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3317 = 6'h35 == _next_can_commit_1_T_1[5:0] ? rob_uop_53_phy_dst : _GEN_3316; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3318 = 6'h36 == _next_can_commit_1_T_1[5:0] ? rob_uop_54_phy_dst : _GEN_3317; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3319 = 6'h37 == _next_can_commit_1_T_1[5:0] ? rob_uop_55_phy_dst : _GEN_3318; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3320 = 6'h38 == _next_can_commit_1_T_1[5:0] ? rob_uop_56_phy_dst : _GEN_3319; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3321 = 6'h39 == _next_can_commit_1_T_1[5:0] ? rob_uop_57_phy_dst : _GEN_3320; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3322 = 6'h3a == _next_can_commit_1_T_1[5:0] ? rob_uop_58_phy_dst : _GEN_3321; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3323 = 6'h3b == _next_can_commit_1_T_1[5:0] ? rob_uop_59_phy_dst : _GEN_3322; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3324 = 6'h3c == _next_can_commit_1_T_1[5:0] ? rob_uop_60_phy_dst : _GEN_3323; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3325 = 6'h3d == _next_can_commit_1_T_1[5:0] ? rob_uop_61_phy_dst : _GEN_3324; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3326 = 6'h3e == _next_can_commit_1_T_1[5:0] ? rob_uop_62_phy_dst : _GEN_3325; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3329 = 6'h1 == _next_can_commit_1_T_1[5:0] ? rob_uop_1_stale_dst : rob_uop_0_stale_dst; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3330 = 6'h2 == _next_can_commit_1_T_1[5:0] ? rob_uop_2_stale_dst : _GEN_3329; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3331 = 6'h3 == _next_can_commit_1_T_1[5:0] ? rob_uop_3_stale_dst : _GEN_3330; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3332 = 6'h4 == _next_can_commit_1_T_1[5:0] ? rob_uop_4_stale_dst : _GEN_3331; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3333 = 6'h5 == _next_can_commit_1_T_1[5:0] ? rob_uop_5_stale_dst : _GEN_3332; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3334 = 6'h6 == _next_can_commit_1_T_1[5:0] ? rob_uop_6_stale_dst : _GEN_3333; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3335 = 6'h7 == _next_can_commit_1_T_1[5:0] ? rob_uop_7_stale_dst : _GEN_3334; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3336 = 6'h8 == _next_can_commit_1_T_1[5:0] ? rob_uop_8_stale_dst : _GEN_3335; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3337 = 6'h9 == _next_can_commit_1_T_1[5:0] ? rob_uop_9_stale_dst : _GEN_3336; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3338 = 6'ha == _next_can_commit_1_T_1[5:0] ? rob_uop_10_stale_dst : _GEN_3337; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3339 = 6'hb == _next_can_commit_1_T_1[5:0] ? rob_uop_11_stale_dst : _GEN_3338; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3340 = 6'hc == _next_can_commit_1_T_1[5:0] ? rob_uop_12_stale_dst : _GEN_3339; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3341 = 6'hd == _next_can_commit_1_T_1[5:0] ? rob_uop_13_stale_dst : _GEN_3340; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3342 = 6'he == _next_can_commit_1_T_1[5:0] ? rob_uop_14_stale_dst : _GEN_3341; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3343 = 6'hf == _next_can_commit_1_T_1[5:0] ? rob_uop_15_stale_dst : _GEN_3342; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3344 = 6'h10 == _next_can_commit_1_T_1[5:0] ? rob_uop_16_stale_dst : _GEN_3343; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3345 = 6'h11 == _next_can_commit_1_T_1[5:0] ? rob_uop_17_stale_dst : _GEN_3344; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3346 = 6'h12 == _next_can_commit_1_T_1[5:0] ? rob_uop_18_stale_dst : _GEN_3345; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3347 = 6'h13 == _next_can_commit_1_T_1[5:0] ? rob_uop_19_stale_dst : _GEN_3346; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3348 = 6'h14 == _next_can_commit_1_T_1[5:0] ? rob_uop_20_stale_dst : _GEN_3347; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3349 = 6'h15 == _next_can_commit_1_T_1[5:0] ? rob_uop_21_stale_dst : _GEN_3348; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3350 = 6'h16 == _next_can_commit_1_T_1[5:0] ? rob_uop_22_stale_dst : _GEN_3349; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3351 = 6'h17 == _next_can_commit_1_T_1[5:0] ? rob_uop_23_stale_dst : _GEN_3350; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3352 = 6'h18 == _next_can_commit_1_T_1[5:0] ? rob_uop_24_stale_dst : _GEN_3351; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3353 = 6'h19 == _next_can_commit_1_T_1[5:0] ? rob_uop_25_stale_dst : _GEN_3352; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3354 = 6'h1a == _next_can_commit_1_T_1[5:0] ? rob_uop_26_stale_dst : _GEN_3353; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3355 = 6'h1b == _next_can_commit_1_T_1[5:0] ? rob_uop_27_stale_dst : _GEN_3354; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3356 = 6'h1c == _next_can_commit_1_T_1[5:0] ? rob_uop_28_stale_dst : _GEN_3355; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3357 = 6'h1d == _next_can_commit_1_T_1[5:0] ? rob_uop_29_stale_dst : _GEN_3356; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3358 = 6'h1e == _next_can_commit_1_T_1[5:0] ? rob_uop_30_stale_dst : _GEN_3357; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3359 = 6'h1f == _next_can_commit_1_T_1[5:0] ? rob_uop_31_stale_dst : _GEN_3358; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3360 = 6'h20 == _next_can_commit_1_T_1[5:0] ? rob_uop_32_stale_dst : _GEN_3359; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3361 = 6'h21 == _next_can_commit_1_T_1[5:0] ? rob_uop_33_stale_dst : _GEN_3360; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3362 = 6'h22 == _next_can_commit_1_T_1[5:0] ? rob_uop_34_stale_dst : _GEN_3361; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3363 = 6'h23 == _next_can_commit_1_T_1[5:0] ? rob_uop_35_stale_dst : _GEN_3362; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3364 = 6'h24 == _next_can_commit_1_T_1[5:0] ? rob_uop_36_stale_dst : _GEN_3363; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3365 = 6'h25 == _next_can_commit_1_T_1[5:0] ? rob_uop_37_stale_dst : _GEN_3364; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3366 = 6'h26 == _next_can_commit_1_T_1[5:0] ? rob_uop_38_stale_dst : _GEN_3365; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3367 = 6'h27 == _next_can_commit_1_T_1[5:0] ? rob_uop_39_stale_dst : _GEN_3366; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3368 = 6'h28 == _next_can_commit_1_T_1[5:0] ? rob_uop_40_stale_dst : _GEN_3367; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3369 = 6'h29 == _next_can_commit_1_T_1[5:0] ? rob_uop_41_stale_dst : _GEN_3368; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3370 = 6'h2a == _next_can_commit_1_T_1[5:0] ? rob_uop_42_stale_dst : _GEN_3369; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3371 = 6'h2b == _next_can_commit_1_T_1[5:0] ? rob_uop_43_stale_dst : _GEN_3370; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3372 = 6'h2c == _next_can_commit_1_T_1[5:0] ? rob_uop_44_stale_dst : _GEN_3371; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3373 = 6'h2d == _next_can_commit_1_T_1[5:0] ? rob_uop_45_stale_dst : _GEN_3372; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3374 = 6'h2e == _next_can_commit_1_T_1[5:0] ? rob_uop_46_stale_dst : _GEN_3373; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3375 = 6'h2f == _next_can_commit_1_T_1[5:0] ? rob_uop_47_stale_dst : _GEN_3374; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3376 = 6'h30 == _next_can_commit_1_T_1[5:0] ? rob_uop_48_stale_dst : _GEN_3375; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3377 = 6'h31 == _next_can_commit_1_T_1[5:0] ? rob_uop_49_stale_dst : _GEN_3376; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3378 = 6'h32 == _next_can_commit_1_T_1[5:0] ? rob_uop_50_stale_dst : _GEN_3377; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3379 = 6'h33 == _next_can_commit_1_T_1[5:0] ? rob_uop_51_stale_dst : _GEN_3378; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3380 = 6'h34 == _next_can_commit_1_T_1[5:0] ? rob_uop_52_stale_dst : _GEN_3379; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3381 = 6'h35 == _next_can_commit_1_T_1[5:0] ? rob_uop_53_stale_dst : _GEN_3380; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3382 = 6'h36 == _next_can_commit_1_T_1[5:0] ? rob_uop_54_stale_dst : _GEN_3381; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3383 = 6'h37 == _next_can_commit_1_T_1[5:0] ? rob_uop_55_stale_dst : _GEN_3382; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3384 = 6'h38 == _next_can_commit_1_T_1[5:0] ? rob_uop_56_stale_dst : _GEN_3383; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3385 = 6'h39 == _next_can_commit_1_T_1[5:0] ? rob_uop_57_stale_dst : _GEN_3384; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3386 = 6'h3a == _next_can_commit_1_T_1[5:0] ? rob_uop_58_stale_dst : _GEN_3385; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3387 = 6'h3b == _next_can_commit_1_T_1[5:0] ? rob_uop_59_stale_dst : _GEN_3386; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3388 = 6'h3c == _next_can_commit_1_T_1[5:0] ? rob_uop_60_stale_dst : _GEN_3387; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3389 = 6'h3d == _next_can_commit_1_T_1[5:0] ? rob_uop_61_stale_dst : _GEN_3388; // @[rob.scala 109:{32,32}]
  wire [6:0] _GEN_3390 = 6'h3e == _next_can_commit_1_T_1[5:0] ? rob_uop_62_stale_dst : _GEN_3389; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3393 = 6'h1 == _next_can_commit_1_T_1[5:0] ? rob_uop_1_arch_dst : rob_uop_0_arch_dst; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3394 = 6'h2 == _next_can_commit_1_T_1[5:0] ? rob_uop_2_arch_dst : _GEN_3393; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3395 = 6'h3 == _next_can_commit_1_T_1[5:0] ? rob_uop_3_arch_dst : _GEN_3394; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3396 = 6'h4 == _next_can_commit_1_T_1[5:0] ? rob_uop_4_arch_dst : _GEN_3395; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3397 = 6'h5 == _next_can_commit_1_T_1[5:0] ? rob_uop_5_arch_dst : _GEN_3396; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3398 = 6'h6 == _next_can_commit_1_T_1[5:0] ? rob_uop_6_arch_dst : _GEN_3397; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3399 = 6'h7 == _next_can_commit_1_T_1[5:0] ? rob_uop_7_arch_dst : _GEN_3398; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3400 = 6'h8 == _next_can_commit_1_T_1[5:0] ? rob_uop_8_arch_dst : _GEN_3399; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3401 = 6'h9 == _next_can_commit_1_T_1[5:0] ? rob_uop_9_arch_dst : _GEN_3400; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3402 = 6'ha == _next_can_commit_1_T_1[5:0] ? rob_uop_10_arch_dst : _GEN_3401; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3403 = 6'hb == _next_can_commit_1_T_1[5:0] ? rob_uop_11_arch_dst : _GEN_3402; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3404 = 6'hc == _next_can_commit_1_T_1[5:0] ? rob_uop_12_arch_dst : _GEN_3403; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3405 = 6'hd == _next_can_commit_1_T_1[5:0] ? rob_uop_13_arch_dst : _GEN_3404; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3406 = 6'he == _next_can_commit_1_T_1[5:0] ? rob_uop_14_arch_dst : _GEN_3405; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3407 = 6'hf == _next_can_commit_1_T_1[5:0] ? rob_uop_15_arch_dst : _GEN_3406; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3408 = 6'h10 == _next_can_commit_1_T_1[5:0] ? rob_uop_16_arch_dst : _GEN_3407; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3409 = 6'h11 == _next_can_commit_1_T_1[5:0] ? rob_uop_17_arch_dst : _GEN_3408; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3410 = 6'h12 == _next_can_commit_1_T_1[5:0] ? rob_uop_18_arch_dst : _GEN_3409; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3411 = 6'h13 == _next_can_commit_1_T_1[5:0] ? rob_uop_19_arch_dst : _GEN_3410; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3412 = 6'h14 == _next_can_commit_1_T_1[5:0] ? rob_uop_20_arch_dst : _GEN_3411; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3413 = 6'h15 == _next_can_commit_1_T_1[5:0] ? rob_uop_21_arch_dst : _GEN_3412; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3414 = 6'h16 == _next_can_commit_1_T_1[5:0] ? rob_uop_22_arch_dst : _GEN_3413; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3415 = 6'h17 == _next_can_commit_1_T_1[5:0] ? rob_uop_23_arch_dst : _GEN_3414; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3416 = 6'h18 == _next_can_commit_1_T_1[5:0] ? rob_uop_24_arch_dst : _GEN_3415; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3417 = 6'h19 == _next_can_commit_1_T_1[5:0] ? rob_uop_25_arch_dst : _GEN_3416; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3418 = 6'h1a == _next_can_commit_1_T_1[5:0] ? rob_uop_26_arch_dst : _GEN_3417; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3419 = 6'h1b == _next_can_commit_1_T_1[5:0] ? rob_uop_27_arch_dst : _GEN_3418; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3420 = 6'h1c == _next_can_commit_1_T_1[5:0] ? rob_uop_28_arch_dst : _GEN_3419; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3421 = 6'h1d == _next_can_commit_1_T_1[5:0] ? rob_uop_29_arch_dst : _GEN_3420; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3422 = 6'h1e == _next_can_commit_1_T_1[5:0] ? rob_uop_30_arch_dst : _GEN_3421; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3423 = 6'h1f == _next_can_commit_1_T_1[5:0] ? rob_uop_31_arch_dst : _GEN_3422; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3424 = 6'h20 == _next_can_commit_1_T_1[5:0] ? rob_uop_32_arch_dst : _GEN_3423; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3425 = 6'h21 == _next_can_commit_1_T_1[5:0] ? rob_uop_33_arch_dst : _GEN_3424; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3426 = 6'h22 == _next_can_commit_1_T_1[5:0] ? rob_uop_34_arch_dst : _GEN_3425; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3427 = 6'h23 == _next_can_commit_1_T_1[5:0] ? rob_uop_35_arch_dst : _GEN_3426; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3428 = 6'h24 == _next_can_commit_1_T_1[5:0] ? rob_uop_36_arch_dst : _GEN_3427; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3429 = 6'h25 == _next_can_commit_1_T_1[5:0] ? rob_uop_37_arch_dst : _GEN_3428; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3430 = 6'h26 == _next_can_commit_1_T_1[5:0] ? rob_uop_38_arch_dst : _GEN_3429; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3431 = 6'h27 == _next_can_commit_1_T_1[5:0] ? rob_uop_39_arch_dst : _GEN_3430; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3432 = 6'h28 == _next_can_commit_1_T_1[5:0] ? rob_uop_40_arch_dst : _GEN_3431; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3433 = 6'h29 == _next_can_commit_1_T_1[5:0] ? rob_uop_41_arch_dst : _GEN_3432; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3434 = 6'h2a == _next_can_commit_1_T_1[5:0] ? rob_uop_42_arch_dst : _GEN_3433; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3435 = 6'h2b == _next_can_commit_1_T_1[5:0] ? rob_uop_43_arch_dst : _GEN_3434; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3436 = 6'h2c == _next_can_commit_1_T_1[5:0] ? rob_uop_44_arch_dst : _GEN_3435; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3437 = 6'h2d == _next_can_commit_1_T_1[5:0] ? rob_uop_45_arch_dst : _GEN_3436; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3438 = 6'h2e == _next_can_commit_1_T_1[5:0] ? rob_uop_46_arch_dst : _GEN_3437; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3439 = 6'h2f == _next_can_commit_1_T_1[5:0] ? rob_uop_47_arch_dst : _GEN_3438; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3440 = 6'h30 == _next_can_commit_1_T_1[5:0] ? rob_uop_48_arch_dst : _GEN_3439; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3441 = 6'h31 == _next_can_commit_1_T_1[5:0] ? rob_uop_49_arch_dst : _GEN_3440; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3442 = 6'h32 == _next_can_commit_1_T_1[5:0] ? rob_uop_50_arch_dst : _GEN_3441; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3443 = 6'h33 == _next_can_commit_1_T_1[5:0] ? rob_uop_51_arch_dst : _GEN_3442; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3444 = 6'h34 == _next_can_commit_1_T_1[5:0] ? rob_uop_52_arch_dst : _GEN_3443; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3445 = 6'h35 == _next_can_commit_1_T_1[5:0] ? rob_uop_53_arch_dst : _GEN_3444; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3446 = 6'h36 == _next_can_commit_1_T_1[5:0] ? rob_uop_54_arch_dst : _GEN_3445; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3447 = 6'h37 == _next_can_commit_1_T_1[5:0] ? rob_uop_55_arch_dst : _GEN_3446; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3448 = 6'h38 == _next_can_commit_1_T_1[5:0] ? rob_uop_56_arch_dst : _GEN_3447; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3449 = 6'h39 == _next_can_commit_1_T_1[5:0] ? rob_uop_57_arch_dst : _GEN_3448; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3450 = 6'h3a == _next_can_commit_1_T_1[5:0] ? rob_uop_58_arch_dst : _GEN_3449; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3451 = 6'h3b == _next_can_commit_1_T_1[5:0] ? rob_uop_59_arch_dst : _GEN_3450; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3452 = 6'h3c == _next_can_commit_1_T_1[5:0] ? rob_uop_60_arch_dst : _GEN_3451; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3453 = 6'h3d == _next_can_commit_1_T_1[5:0] ? rob_uop_61_arch_dst : _GEN_3452; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_3454 = 6'h3e == _next_can_commit_1_T_1[5:0] ? rob_uop_62_arch_dst : _GEN_3453; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4097 = 6'h1 == _next_can_commit_1_T_1[5:0] ? rob_uop_1_dst_value : rob_uop_0_dst_value; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4098 = 6'h2 == _next_can_commit_1_T_1[5:0] ? rob_uop_2_dst_value : _GEN_4097; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4099 = 6'h3 == _next_can_commit_1_T_1[5:0] ? rob_uop_3_dst_value : _GEN_4098; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4100 = 6'h4 == _next_can_commit_1_T_1[5:0] ? rob_uop_4_dst_value : _GEN_4099; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4101 = 6'h5 == _next_can_commit_1_T_1[5:0] ? rob_uop_5_dst_value : _GEN_4100; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4102 = 6'h6 == _next_can_commit_1_T_1[5:0] ? rob_uop_6_dst_value : _GEN_4101; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4103 = 6'h7 == _next_can_commit_1_T_1[5:0] ? rob_uop_7_dst_value : _GEN_4102; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4104 = 6'h8 == _next_can_commit_1_T_1[5:0] ? rob_uop_8_dst_value : _GEN_4103; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4105 = 6'h9 == _next_can_commit_1_T_1[5:0] ? rob_uop_9_dst_value : _GEN_4104; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4106 = 6'ha == _next_can_commit_1_T_1[5:0] ? rob_uop_10_dst_value : _GEN_4105; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4107 = 6'hb == _next_can_commit_1_T_1[5:0] ? rob_uop_11_dst_value : _GEN_4106; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4108 = 6'hc == _next_can_commit_1_T_1[5:0] ? rob_uop_12_dst_value : _GEN_4107; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4109 = 6'hd == _next_can_commit_1_T_1[5:0] ? rob_uop_13_dst_value : _GEN_4108; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4110 = 6'he == _next_can_commit_1_T_1[5:0] ? rob_uop_14_dst_value : _GEN_4109; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4111 = 6'hf == _next_can_commit_1_T_1[5:0] ? rob_uop_15_dst_value : _GEN_4110; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4112 = 6'h10 == _next_can_commit_1_T_1[5:0] ? rob_uop_16_dst_value : _GEN_4111; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4113 = 6'h11 == _next_can_commit_1_T_1[5:0] ? rob_uop_17_dst_value : _GEN_4112; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4114 = 6'h12 == _next_can_commit_1_T_1[5:0] ? rob_uop_18_dst_value : _GEN_4113; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4115 = 6'h13 == _next_can_commit_1_T_1[5:0] ? rob_uop_19_dst_value : _GEN_4114; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4116 = 6'h14 == _next_can_commit_1_T_1[5:0] ? rob_uop_20_dst_value : _GEN_4115; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4117 = 6'h15 == _next_can_commit_1_T_1[5:0] ? rob_uop_21_dst_value : _GEN_4116; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4118 = 6'h16 == _next_can_commit_1_T_1[5:0] ? rob_uop_22_dst_value : _GEN_4117; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4119 = 6'h17 == _next_can_commit_1_T_1[5:0] ? rob_uop_23_dst_value : _GEN_4118; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4120 = 6'h18 == _next_can_commit_1_T_1[5:0] ? rob_uop_24_dst_value : _GEN_4119; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4121 = 6'h19 == _next_can_commit_1_T_1[5:0] ? rob_uop_25_dst_value : _GEN_4120; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4122 = 6'h1a == _next_can_commit_1_T_1[5:0] ? rob_uop_26_dst_value : _GEN_4121; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4123 = 6'h1b == _next_can_commit_1_T_1[5:0] ? rob_uop_27_dst_value : _GEN_4122; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4124 = 6'h1c == _next_can_commit_1_T_1[5:0] ? rob_uop_28_dst_value : _GEN_4123; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4125 = 6'h1d == _next_can_commit_1_T_1[5:0] ? rob_uop_29_dst_value : _GEN_4124; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4126 = 6'h1e == _next_can_commit_1_T_1[5:0] ? rob_uop_30_dst_value : _GEN_4125; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4127 = 6'h1f == _next_can_commit_1_T_1[5:0] ? rob_uop_31_dst_value : _GEN_4126; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4128 = 6'h20 == _next_can_commit_1_T_1[5:0] ? rob_uop_32_dst_value : _GEN_4127; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4129 = 6'h21 == _next_can_commit_1_T_1[5:0] ? rob_uop_33_dst_value : _GEN_4128; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4130 = 6'h22 == _next_can_commit_1_T_1[5:0] ? rob_uop_34_dst_value : _GEN_4129; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4131 = 6'h23 == _next_can_commit_1_T_1[5:0] ? rob_uop_35_dst_value : _GEN_4130; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4132 = 6'h24 == _next_can_commit_1_T_1[5:0] ? rob_uop_36_dst_value : _GEN_4131; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4133 = 6'h25 == _next_can_commit_1_T_1[5:0] ? rob_uop_37_dst_value : _GEN_4132; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4134 = 6'h26 == _next_can_commit_1_T_1[5:0] ? rob_uop_38_dst_value : _GEN_4133; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4135 = 6'h27 == _next_can_commit_1_T_1[5:0] ? rob_uop_39_dst_value : _GEN_4134; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4136 = 6'h28 == _next_can_commit_1_T_1[5:0] ? rob_uop_40_dst_value : _GEN_4135; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4137 = 6'h29 == _next_can_commit_1_T_1[5:0] ? rob_uop_41_dst_value : _GEN_4136; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4138 = 6'h2a == _next_can_commit_1_T_1[5:0] ? rob_uop_42_dst_value : _GEN_4137; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4139 = 6'h2b == _next_can_commit_1_T_1[5:0] ? rob_uop_43_dst_value : _GEN_4138; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4140 = 6'h2c == _next_can_commit_1_T_1[5:0] ? rob_uop_44_dst_value : _GEN_4139; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4141 = 6'h2d == _next_can_commit_1_T_1[5:0] ? rob_uop_45_dst_value : _GEN_4140; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4142 = 6'h2e == _next_can_commit_1_T_1[5:0] ? rob_uop_46_dst_value : _GEN_4141; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4143 = 6'h2f == _next_can_commit_1_T_1[5:0] ? rob_uop_47_dst_value : _GEN_4142; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4144 = 6'h30 == _next_can_commit_1_T_1[5:0] ? rob_uop_48_dst_value : _GEN_4143; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4145 = 6'h31 == _next_can_commit_1_T_1[5:0] ? rob_uop_49_dst_value : _GEN_4144; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4146 = 6'h32 == _next_can_commit_1_T_1[5:0] ? rob_uop_50_dst_value : _GEN_4145; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4147 = 6'h33 == _next_can_commit_1_T_1[5:0] ? rob_uop_51_dst_value : _GEN_4146; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4148 = 6'h34 == _next_can_commit_1_T_1[5:0] ? rob_uop_52_dst_value : _GEN_4147; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4149 = 6'h35 == _next_can_commit_1_T_1[5:0] ? rob_uop_53_dst_value : _GEN_4148; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4150 = 6'h36 == _next_can_commit_1_T_1[5:0] ? rob_uop_54_dst_value : _GEN_4149; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4151 = 6'h37 == _next_can_commit_1_T_1[5:0] ? rob_uop_55_dst_value : _GEN_4150; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4152 = 6'h38 == _next_can_commit_1_T_1[5:0] ? rob_uop_56_dst_value : _GEN_4151; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4153 = 6'h39 == _next_can_commit_1_T_1[5:0] ? rob_uop_57_dst_value : _GEN_4152; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4154 = 6'h3a == _next_can_commit_1_T_1[5:0] ? rob_uop_58_dst_value : _GEN_4153; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4155 = 6'h3b == _next_can_commit_1_T_1[5:0] ? rob_uop_59_dst_value : _GEN_4154; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4156 = 6'h3c == _next_can_commit_1_T_1[5:0] ? rob_uop_60_dst_value : _GEN_4155; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4157 = 6'h3d == _next_can_commit_1_T_1[5:0] ? rob_uop_61_dst_value : _GEN_4156; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4158 = 6'h3e == _next_can_commit_1_T_1[5:0] ? rob_uop_62_dst_value : _GEN_4157; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4161 = 6'h1 == _next_can_commit_1_T_1[5:0] ? rob_uop_1_src1_value : rob_uop_0_src1_value; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4162 = 6'h2 == _next_can_commit_1_T_1[5:0] ? rob_uop_2_src1_value : _GEN_4161; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4163 = 6'h3 == _next_can_commit_1_T_1[5:0] ? rob_uop_3_src1_value : _GEN_4162; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4164 = 6'h4 == _next_can_commit_1_T_1[5:0] ? rob_uop_4_src1_value : _GEN_4163; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4165 = 6'h5 == _next_can_commit_1_T_1[5:0] ? rob_uop_5_src1_value : _GEN_4164; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4166 = 6'h6 == _next_can_commit_1_T_1[5:0] ? rob_uop_6_src1_value : _GEN_4165; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4167 = 6'h7 == _next_can_commit_1_T_1[5:0] ? rob_uop_7_src1_value : _GEN_4166; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4168 = 6'h8 == _next_can_commit_1_T_1[5:0] ? rob_uop_8_src1_value : _GEN_4167; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4169 = 6'h9 == _next_can_commit_1_T_1[5:0] ? rob_uop_9_src1_value : _GEN_4168; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4170 = 6'ha == _next_can_commit_1_T_1[5:0] ? rob_uop_10_src1_value : _GEN_4169; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4171 = 6'hb == _next_can_commit_1_T_1[5:0] ? rob_uop_11_src1_value : _GEN_4170; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4172 = 6'hc == _next_can_commit_1_T_1[5:0] ? rob_uop_12_src1_value : _GEN_4171; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4173 = 6'hd == _next_can_commit_1_T_1[5:0] ? rob_uop_13_src1_value : _GEN_4172; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4174 = 6'he == _next_can_commit_1_T_1[5:0] ? rob_uop_14_src1_value : _GEN_4173; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4175 = 6'hf == _next_can_commit_1_T_1[5:0] ? rob_uop_15_src1_value : _GEN_4174; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4176 = 6'h10 == _next_can_commit_1_T_1[5:0] ? rob_uop_16_src1_value : _GEN_4175; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4177 = 6'h11 == _next_can_commit_1_T_1[5:0] ? rob_uop_17_src1_value : _GEN_4176; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4178 = 6'h12 == _next_can_commit_1_T_1[5:0] ? rob_uop_18_src1_value : _GEN_4177; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4179 = 6'h13 == _next_can_commit_1_T_1[5:0] ? rob_uop_19_src1_value : _GEN_4178; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4180 = 6'h14 == _next_can_commit_1_T_1[5:0] ? rob_uop_20_src1_value : _GEN_4179; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4181 = 6'h15 == _next_can_commit_1_T_1[5:0] ? rob_uop_21_src1_value : _GEN_4180; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4182 = 6'h16 == _next_can_commit_1_T_1[5:0] ? rob_uop_22_src1_value : _GEN_4181; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4183 = 6'h17 == _next_can_commit_1_T_1[5:0] ? rob_uop_23_src1_value : _GEN_4182; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4184 = 6'h18 == _next_can_commit_1_T_1[5:0] ? rob_uop_24_src1_value : _GEN_4183; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4185 = 6'h19 == _next_can_commit_1_T_1[5:0] ? rob_uop_25_src1_value : _GEN_4184; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4186 = 6'h1a == _next_can_commit_1_T_1[5:0] ? rob_uop_26_src1_value : _GEN_4185; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4187 = 6'h1b == _next_can_commit_1_T_1[5:0] ? rob_uop_27_src1_value : _GEN_4186; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4188 = 6'h1c == _next_can_commit_1_T_1[5:0] ? rob_uop_28_src1_value : _GEN_4187; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4189 = 6'h1d == _next_can_commit_1_T_1[5:0] ? rob_uop_29_src1_value : _GEN_4188; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4190 = 6'h1e == _next_can_commit_1_T_1[5:0] ? rob_uop_30_src1_value : _GEN_4189; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4191 = 6'h1f == _next_can_commit_1_T_1[5:0] ? rob_uop_31_src1_value : _GEN_4190; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4192 = 6'h20 == _next_can_commit_1_T_1[5:0] ? rob_uop_32_src1_value : _GEN_4191; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4193 = 6'h21 == _next_can_commit_1_T_1[5:0] ? rob_uop_33_src1_value : _GEN_4192; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4194 = 6'h22 == _next_can_commit_1_T_1[5:0] ? rob_uop_34_src1_value : _GEN_4193; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4195 = 6'h23 == _next_can_commit_1_T_1[5:0] ? rob_uop_35_src1_value : _GEN_4194; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4196 = 6'h24 == _next_can_commit_1_T_1[5:0] ? rob_uop_36_src1_value : _GEN_4195; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4197 = 6'h25 == _next_can_commit_1_T_1[5:0] ? rob_uop_37_src1_value : _GEN_4196; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4198 = 6'h26 == _next_can_commit_1_T_1[5:0] ? rob_uop_38_src1_value : _GEN_4197; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4199 = 6'h27 == _next_can_commit_1_T_1[5:0] ? rob_uop_39_src1_value : _GEN_4198; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4200 = 6'h28 == _next_can_commit_1_T_1[5:0] ? rob_uop_40_src1_value : _GEN_4199; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4201 = 6'h29 == _next_can_commit_1_T_1[5:0] ? rob_uop_41_src1_value : _GEN_4200; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4202 = 6'h2a == _next_can_commit_1_T_1[5:0] ? rob_uop_42_src1_value : _GEN_4201; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4203 = 6'h2b == _next_can_commit_1_T_1[5:0] ? rob_uop_43_src1_value : _GEN_4202; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4204 = 6'h2c == _next_can_commit_1_T_1[5:0] ? rob_uop_44_src1_value : _GEN_4203; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4205 = 6'h2d == _next_can_commit_1_T_1[5:0] ? rob_uop_45_src1_value : _GEN_4204; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4206 = 6'h2e == _next_can_commit_1_T_1[5:0] ? rob_uop_46_src1_value : _GEN_4205; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4207 = 6'h2f == _next_can_commit_1_T_1[5:0] ? rob_uop_47_src1_value : _GEN_4206; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4208 = 6'h30 == _next_can_commit_1_T_1[5:0] ? rob_uop_48_src1_value : _GEN_4207; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4209 = 6'h31 == _next_can_commit_1_T_1[5:0] ? rob_uop_49_src1_value : _GEN_4208; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4210 = 6'h32 == _next_can_commit_1_T_1[5:0] ? rob_uop_50_src1_value : _GEN_4209; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4211 = 6'h33 == _next_can_commit_1_T_1[5:0] ? rob_uop_51_src1_value : _GEN_4210; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4212 = 6'h34 == _next_can_commit_1_T_1[5:0] ? rob_uop_52_src1_value : _GEN_4211; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4213 = 6'h35 == _next_can_commit_1_T_1[5:0] ? rob_uop_53_src1_value : _GEN_4212; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4214 = 6'h36 == _next_can_commit_1_T_1[5:0] ? rob_uop_54_src1_value : _GEN_4213; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4215 = 6'h37 == _next_can_commit_1_T_1[5:0] ? rob_uop_55_src1_value : _GEN_4214; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4216 = 6'h38 == _next_can_commit_1_T_1[5:0] ? rob_uop_56_src1_value : _GEN_4215; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4217 = 6'h39 == _next_can_commit_1_T_1[5:0] ? rob_uop_57_src1_value : _GEN_4216; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4218 = 6'h3a == _next_can_commit_1_T_1[5:0] ? rob_uop_58_src1_value : _GEN_4217; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4219 = 6'h3b == _next_can_commit_1_T_1[5:0] ? rob_uop_59_src1_value : _GEN_4218; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4220 = 6'h3c == _next_can_commit_1_T_1[5:0] ? rob_uop_60_src1_value : _GEN_4219; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4221 = 6'h3d == _next_can_commit_1_T_1[5:0] ? rob_uop_61_src1_value : _GEN_4220; // @[rob.scala 109:{32,32}]
  wire [63:0] _GEN_4222 = 6'h3e == _next_can_commit_1_T_1[5:0] ? rob_uop_62_src1_value : _GEN_4221; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4481 = 6'h1 == _next_can_commit_1_T_1[5:0] ? rob_uop_1_alu_sel : rob_uop_0_alu_sel; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4482 = 6'h2 == _next_can_commit_1_T_1[5:0] ? rob_uop_2_alu_sel : _GEN_4481; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4483 = 6'h3 == _next_can_commit_1_T_1[5:0] ? rob_uop_3_alu_sel : _GEN_4482; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4484 = 6'h4 == _next_can_commit_1_T_1[5:0] ? rob_uop_4_alu_sel : _GEN_4483; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4485 = 6'h5 == _next_can_commit_1_T_1[5:0] ? rob_uop_5_alu_sel : _GEN_4484; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4486 = 6'h6 == _next_can_commit_1_T_1[5:0] ? rob_uop_6_alu_sel : _GEN_4485; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4487 = 6'h7 == _next_can_commit_1_T_1[5:0] ? rob_uop_7_alu_sel : _GEN_4486; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4488 = 6'h8 == _next_can_commit_1_T_1[5:0] ? rob_uop_8_alu_sel : _GEN_4487; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4489 = 6'h9 == _next_can_commit_1_T_1[5:0] ? rob_uop_9_alu_sel : _GEN_4488; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4490 = 6'ha == _next_can_commit_1_T_1[5:0] ? rob_uop_10_alu_sel : _GEN_4489; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4491 = 6'hb == _next_can_commit_1_T_1[5:0] ? rob_uop_11_alu_sel : _GEN_4490; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4492 = 6'hc == _next_can_commit_1_T_1[5:0] ? rob_uop_12_alu_sel : _GEN_4491; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4493 = 6'hd == _next_can_commit_1_T_1[5:0] ? rob_uop_13_alu_sel : _GEN_4492; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4494 = 6'he == _next_can_commit_1_T_1[5:0] ? rob_uop_14_alu_sel : _GEN_4493; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4495 = 6'hf == _next_can_commit_1_T_1[5:0] ? rob_uop_15_alu_sel : _GEN_4494; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4496 = 6'h10 == _next_can_commit_1_T_1[5:0] ? rob_uop_16_alu_sel : _GEN_4495; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4497 = 6'h11 == _next_can_commit_1_T_1[5:0] ? rob_uop_17_alu_sel : _GEN_4496; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4498 = 6'h12 == _next_can_commit_1_T_1[5:0] ? rob_uop_18_alu_sel : _GEN_4497; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4499 = 6'h13 == _next_can_commit_1_T_1[5:0] ? rob_uop_19_alu_sel : _GEN_4498; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4500 = 6'h14 == _next_can_commit_1_T_1[5:0] ? rob_uop_20_alu_sel : _GEN_4499; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4501 = 6'h15 == _next_can_commit_1_T_1[5:0] ? rob_uop_21_alu_sel : _GEN_4500; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4502 = 6'h16 == _next_can_commit_1_T_1[5:0] ? rob_uop_22_alu_sel : _GEN_4501; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4503 = 6'h17 == _next_can_commit_1_T_1[5:0] ? rob_uop_23_alu_sel : _GEN_4502; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4504 = 6'h18 == _next_can_commit_1_T_1[5:0] ? rob_uop_24_alu_sel : _GEN_4503; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4505 = 6'h19 == _next_can_commit_1_T_1[5:0] ? rob_uop_25_alu_sel : _GEN_4504; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4506 = 6'h1a == _next_can_commit_1_T_1[5:0] ? rob_uop_26_alu_sel : _GEN_4505; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4507 = 6'h1b == _next_can_commit_1_T_1[5:0] ? rob_uop_27_alu_sel : _GEN_4506; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4508 = 6'h1c == _next_can_commit_1_T_1[5:0] ? rob_uop_28_alu_sel : _GEN_4507; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4509 = 6'h1d == _next_can_commit_1_T_1[5:0] ? rob_uop_29_alu_sel : _GEN_4508; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4510 = 6'h1e == _next_can_commit_1_T_1[5:0] ? rob_uop_30_alu_sel : _GEN_4509; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4511 = 6'h1f == _next_can_commit_1_T_1[5:0] ? rob_uop_31_alu_sel : _GEN_4510; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4512 = 6'h20 == _next_can_commit_1_T_1[5:0] ? rob_uop_32_alu_sel : _GEN_4511; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4513 = 6'h21 == _next_can_commit_1_T_1[5:0] ? rob_uop_33_alu_sel : _GEN_4512; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4514 = 6'h22 == _next_can_commit_1_T_1[5:0] ? rob_uop_34_alu_sel : _GEN_4513; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4515 = 6'h23 == _next_can_commit_1_T_1[5:0] ? rob_uop_35_alu_sel : _GEN_4514; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4516 = 6'h24 == _next_can_commit_1_T_1[5:0] ? rob_uop_36_alu_sel : _GEN_4515; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4517 = 6'h25 == _next_can_commit_1_T_1[5:0] ? rob_uop_37_alu_sel : _GEN_4516; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4518 = 6'h26 == _next_can_commit_1_T_1[5:0] ? rob_uop_38_alu_sel : _GEN_4517; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4519 = 6'h27 == _next_can_commit_1_T_1[5:0] ? rob_uop_39_alu_sel : _GEN_4518; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4520 = 6'h28 == _next_can_commit_1_T_1[5:0] ? rob_uop_40_alu_sel : _GEN_4519; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4521 = 6'h29 == _next_can_commit_1_T_1[5:0] ? rob_uop_41_alu_sel : _GEN_4520; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4522 = 6'h2a == _next_can_commit_1_T_1[5:0] ? rob_uop_42_alu_sel : _GEN_4521; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4523 = 6'h2b == _next_can_commit_1_T_1[5:0] ? rob_uop_43_alu_sel : _GEN_4522; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4524 = 6'h2c == _next_can_commit_1_T_1[5:0] ? rob_uop_44_alu_sel : _GEN_4523; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4525 = 6'h2d == _next_can_commit_1_T_1[5:0] ? rob_uop_45_alu_sel : _GEN_4524; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4526 = 6'h2e == _next_can_commit_1_T_1[5:0] ? rob_uop_46_alu_sel : _GEN_4525; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4527 = 6'h2f == _next_can_commit_1_T_1[5:0] ? rob_uop_47_alu_sel : _GEN_4526; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4528 = 6'h30 == _next_can_commit_1_T_1[5:0] ? rob_uop_48_alu_sel : _GEN_4527; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4529 = 6'h31 == _next_can_commit_1_T_1[5:0] ? rob_uop_49_alu_sel : _GEN_4528; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4530 = 6'h32 == _next_can_commit_1_T_1[5:0] ? rob_uop_50_alu_sel : _GEN_4529; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4531 = 6'h33 == _next_can_commit_1_T_1[5:0] ? rob_uop_51_alu_sel : _GEN_4530; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4532 = 6'h34 == _next_can_commit_1_T_1[5:0] ? rob_uop_52_alu_sel : _GEN_4531; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4533 = 6'h35 == _next_can_commit_1_T_1[5:0] ? rob_uop_53_alu_sel : _GEN_4532; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4534 = 6'h36 == _next_can_commit_1_T_1[5:0] ? rob_uop_54_alu_sel : _GEN_4533; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4535 = 6'h37 == _next_can_commit_1_T_1[5:0] ? rob_uop_55_alu_sel : _GEN_4534; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4536 = 6'h38 == _next_can_commit_1_T_1[5:0] ? rob_uop_56_alu_sel : _GEN_4535; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4537 = 6'h39 == _next_can_commit_1_T_1[5:0] ? rob_uop_57_alu_sel : _GEN_4536; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4538 = 6'h3a == _next_can_commit_1_T_1[5:0] ? rob_uop_58_alu_sel : _GEN_4537; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4539 = 6'h3b == _next_can_commit_1_T_1[5:0] ? rob_uop_59_alu_sel : _GEN_4538; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4540 = 6'h3c == _next_can_commit_1_T_1[5:0] ? rob_uop_60_alu_sel : _GEN_4539; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4541 = 6'h3d == _next_can_commit_1_T_1[5:0] ? rob_uop_61_alu_sel : _GEN_4540; // @[rob.scala 109:{32,32}]
  wire [4:0] _GEN_4542 = 6'h3e == _next_can_commit_1_T_1[5:0] ? rob_uop_62_alu_sel : _GEN_4541; // @[rob.scala 109:{32,32}]
  wire [6:0] this_num_to_roll_back = {{5'd0}, _this_num_to_roll_back_T_17}; // @[rob.scala 66:37 73:27]
  wire [6:0] _GEN_5249 = 6'h1 == _next_rob_state_T_10[5:0] ? rob_uop_1_phy_dst : rob_uop_0_phy_dst; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5250 = 6'h2 == _next_rob_state_T_10[5:0] ? rob_uop_2_phy_dst : _GEN_5249; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5251 = 6'h3 == _next_rob_state_T_10[5:0] ? rob_uop_3_phy_dst : _GEN_5250; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5252 = 6'h4 == _next_rob_state_T_10[5:0] ? rob_uop_4_phy_dst : _GEN_5251; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5253 = 6'h5 == _next_rob_state_T_10[5:0] ? rob_uop_5_phy_dst : _GEN_5252; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5254 = 6'h6 == _next_rob_state_T_10[5:0] ? rob_uop_6_phy_dst : _GEN_5253; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5255 = 6'h7 == _next_rob_state_T_10[5:0] ? rob_uop_7_phy_dst : _GEN_5254; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5256 = 6'h8 == _next_rob_state_T_10[5:0] ? rob_uop_8_phy_dst : _GEN_5255; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5257 = 6'h9 == _next_rob_state_T_10[5:0] ? rob_uop_9_phy_dst : _GEN_5256; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5258 = 6'ha == _next_rob_state_T_10[5:0] ? rob_uop_10_phy_dst : _GEN_5257; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5259 = 6'hb == _next_rob_state_T_10[5:0] ? rob_uop_11_phy_dst : _GEN_5258; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5260 = 6'hc == _next_rob_state_T_10[5:0] ? rob_uop_12_phy_dst : _GEN_5259; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5261 = 6'hd == _next_rob_state_T_10[5:0] ? rob_uop_13_phy_dst : _GEN_5260; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5262 = 6'he == _next_rob_state_T_10[5:0] ? rob_uop_14_phy_dst : _GEN_5261; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5263 = 6'hf == _next_rob_state_T_10[5:0] ? rob_uop_15_phy_dst : _GEN_5262; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5264 = 6'h10 == _next_rob_state_T_10[5:0] ? rob_uop_16_phy_dst : _GEN_5263; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5265 = 6'h11 == _next_rob_state_T_10[5:0] ? rob_uop_17_phy_dst : _GEN_5264; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5266 = 6'h12 == _next_rob_state_T_10[5:0] ? rob_uop_18_phy_dst : _GEN_5265; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5267 = 6'h13 == _next_rob_state_T_10[5:0] ? rob_uop_19_phy_dst : _GEN_5266; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5268 = 6'h14 == _next_rob_state_T_10[5:0] ? rob_uop_20_phy_dst : _GEN_5267; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5269 = 6'h15 == _next_rob_state_T_10[5:0] ? rob_uop_21_phy_dst : _GEN_5268; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5270 = 6'h16 == _next_rob_state_T_10[5:0] ? rob_uop_22_phy_dst : _GEN_5269; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5271 = 6'h17 == _next_rob_state_T_10[5:0] ? rob_uop_23_phy_dst : _GEN_5270; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5272 = 6'h18 == _next_rob_state_T_10[5:0] ? rob_uop_24_phy_dst : _GEN_5271; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5273 = 6'h19 == _next_rob_state_T_10[5:0] ? rob_uop_25_phy_dst : _GEN_5272; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5274 = 6'h1a == _next_rob_state_T_10[5:0] ? rob_uop_26_phy_dst : _GEN_5273; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5275 = 6'h1b == _next_rob_state_T_10[5:0] ? rob_uop_27_phy_dst : _GEN_5274; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5276 = 6'h1c == _next_rob_state_T_10[5:0] ? rob_uop_28_phy_dst : _GEN_5275; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5277 = 6'h1d == _next_rob_state_T_10[5:0] ? rob_uop_29_phy_dst : _GEN_5276; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5278 = 6'h1e == _next_rob_state_T_10[5:0] ? rob_uop_30_phy_dst : _GEN_5277; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5279 = 6'h1f == _next_rob_state_T_10[5:0] ? rob_uop_31_phy_dst : _GEN_5278; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5280 = 6'h20 == _next_rob_state_T_10[5:0] ? rob_uop_32_phy_dst : _GEN_5279; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5281 = 6'h21 == _next_rob_state_T_10[5:0] ? rob_uop_33_phy_dst : _GEN_5280; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5282 = 6'h22 == _next_rob_state_T_10[5:0] ? rob_uop_34_phy_dst : _GEN_5281; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5283 = 6'h23 == _next_rob_state_T_10[5:0] ? rob_uop_35_phy_dst : _GEN_5282; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5284 = 6'h24 == _next_rob_state_T_10[5:0] ? rob_uop_36_phy_dst : _GEN_5283; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5285 = 6'h25 == _next_rob_state_T_10[5:0] ? rob_uop_37_phy_dst : _GEN_5284; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5286 = 6'h26 == _next_rob_state_T_10[5:0] ? rob_uop_38_phy_dst : _GEN_5285; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5287 = 6'h27 == _next_rob_state_T_10[5:0] ? rob_uop_39_phy_dst : _GEN_5286; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5288 = 6'h28 == _next_rob_state_T_10[5:0] ? rob_uop_40_phy_dst : _GEN_5287; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5289 = 6'h29 == _next_rob_state_T_10[5:0] ? rob_uop_41_phy_dst : _GEN_5288; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5290 = 6'h2a == _next_rob_state_T_10[5:0] ? rob_uop_42_phy_dst : _GEN_5289; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5291 = 6'h2b == _next_rob_state_T_10[5:0] ? rob_uop_43_phy_dst : _GEN_5290; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5292 = 6'h2c == _next_rob_state_T_10[5:0] ? rob_uop_44_phy_dst : _GEN_5291; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5293 = 6'h2d == _next_rob_state_T_10[5:0] ? rob_uop_45_phy_dst : _GEN_5292; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5294 = 6'h2e == _next_rob_state_T_10[5:0] ? rob_uop_46_phy_dst : _GEN_5293; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5295 = 6'h2f == _next_rob_state_T_10[5:0] ? rob_uop_47_phy_dst : _GEN_5294; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5296 = 6'h30 == _next_rob_state_T_10[5:0] ? rob_uop_48_phy_dst : _GEN_5295; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5297 = 6'h31 == _next_rob_state_T_10[5:0] ? rob_uop_49_phy_dst : _GEN_5296; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5298 = 6'h32 == _next_rob_state_T_10[5:0] ? rob_uop_50_phy_dst : _GEN_5297; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5299 = 6'h33 == _next_rob_state_T_10[5:0] ? rob_uop_51_phy_dst : _GEN_5298; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5300 = 6'h34 == _next_rob_state_T_10[5:0] ? rob_uop_52_phy_dst : _GEN_5299; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5301 = 6'h35 == _next_rob_state_T_10[5:0] ? rob_uop_53_phy_dst : _GEN_5300; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5302 = 6'h36 == _next_rob_state_T_10[5:0] ? rob_uop_54_phy_dst : _GEN_5301; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5303 = 6'h37 == _next_rob_state_T_10[5:0] ? rob_uop_55_phy_dst : _GEN_5302; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5304 = 6'h38 == _next_rob_state_T_10[5:0] ? rob_uop_56_phy_dst : _GEN_5303; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5305 = 6'h39 == _next_rob_state_T_10[5:0] ? rob_uop_57_phy_dst : _GEN_5304; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5306 = 6'h3a == _next_rob_state_T_10[5:0] ? rob_uop_58_phy_dst : _GEN_5305; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5307 = 6'h3b == _next_rob_state_T_10[5:0] ? rob_uop_59_phy_dst : _GEN_5306; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5308 = 6'h3c == _next_rob_state_T_10[5:0] ? rob_uop_60_phy_dst : _GEN_5307; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5309 = 6'h3d == _next_rob_state_T_10[5:0] ? rob_uop_61_phy_dst : _GEN_5308; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5310 = 6'h3e == _next_rob_state_T_10[5:0] ? rob_uop_62_phy_dst : _GEN_5309; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5313 = 6'h1 == _next_rob_state_T_10[5:0] ? rob_uop_1_stale_dst : rob_uop_0_stale_dst; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5314 = 6'h2 == _next_rob_state_T_10[5:0] ? rob_uop_2_stale_dst : _GEN_5313; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5315 = 6'h3 == _next_rob_state_T_10[5:0] ? rob_uop_3_stale_dst : _GEN_5314; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5316 = 6'h4 == _next_rob_state_T_10[5:0] ? rob_uop_4_stale_dst : _GEN_5315; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5317 = 6'h5 == _next_rob_state_T_10[5:0] ? rob_uop_5_stale_dst : _GEN_5316; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5318 = 6'h6 == _next_rob_state_T_10[5:0] ? rob_uop_6_stale_dst : _GEN_5317; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5319 = 6'h7 == _next_rob_state_T_10[5:0] ? rob_uop_7_stale_dst : _GEN_5318; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5320 = 6'h8 == _next_rob_state_T_10[5:0] ? rob_uop_8_stale_dst : _GEN_5319; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5321 = 6'h9 == _next_rob_state_T_10[5:0] ? rob_uop_9_stale_dst : _GEN_5320; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5322 = 6'ha == _next_rob_state_T_10[5:0] ? rob_uop_10_stale_dst : _GEN_5321; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5323 = 6'hb == _next_rob_state_T_10[5:0] ? rob_uop_11_stale_dst : _GEN_5322; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5324 = 6'hc == _next_rob_state_T_10[5:0] ? rob_uop_12_stale_dst : _GEN_5323; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5325 = 6'hd == _next_rob_state_T_10[5:0] ? rob_uop_13_stale_dst : _GEN_5324; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5326 = 6'he == _next_rob_state_T_10[5:0] ? rob_uop_14_stale_dst : _GEN_5325; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5327 = 6'hf == _next_rob_state_T_10[5:0] ? rob_uop_15_stale_dst : _GEN_5326; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5328 = 6'h10 == _next_rob_state_T_10[5:0] ? rob_uop_16_stale_dst : _GEN_5327; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5329 = 6'h11 == _next_rob_state_T_10[5:0] ? rob_uop_17_stale_dst : _GEN_5328; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5330 = 6'h12 == _next_rob_state_T_10[5:0] ? rob_uop_18_stale_dst : _GEN_5329; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5331 = 6'h13 == _next_rob_state_T_10[5:0] ? rob_uop_19_stale_dst : _GEN_5330; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5332 = 6'h14 == _next_rob_state_T_10[5:0] ? rob_uop_20_stale_dst : _GEN_5331; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5333 = 6'h15 == _next_rob_state_T_10[5:0] ? rob_uop_21_stale_dst : _GEN_5332; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5334 = 6'h16 == _next_rob_state_T_10[5:0] ? rob_uop_22_stale_dst : _GEN_5333; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5335 = 6'h17 == _next_rob_state_T_10[5:0] ? rob_uop_23_stale_dst : _GEN_5334; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5336 = 6'h18 == _next_rob_state_T_10[5:0] ? rob_uop_24_stale_dst : _GEN_5335; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5337 = 6'h19 == _next_rob_state_T_10[5:0] ? rob_uop_25_stale_dst : _GEN_5336; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5338 = 6'h1a == _next_rob_state_T_10[5:0] ? rob_uop_26_stale_dst : _GEN_5337; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5339 = 6'h1b == _next_rob_state_T_10[5:0] ? rob_uop_27_stale_dst : _GEN_5338; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5340 = 6'h1c == _next_rob_state_T_10[5:0] ? rob_uop_28_stale_dst : _GEN_5339; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5341 = 6'h1d == _next_rob_state_T_10[5:0] ? rob_uop_29_stale_dst : _GEN_5340; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5342 = 6'h1e == _next_rob_state_T_10[5:0] ? rob_uop_30_stale_dst : _GEN_5341; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5343 = 6'h1f == _next_rob_state_T_10[5:0] ? rob_uop_31_stale_dst : _GEN_5342; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5344 = 6'h20 == _next_rob_state_T_10[5:0] ? rob_uop_32_stale_dst : _GEN_5343; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5345 = 6'h21 == _next_rob_state_T_10[5:0] ? rob_uop_33_stale_dst : _GEN_5344; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5346 = 6'h22 == _next_rob_state_T_10[5:0] ? rob_uop_34_stale_dst : _GEN_5345; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5347 = 6'h23 == _next_rob_state_T_10[5:0] ? rob_uop_35_stale_dst : _GEN_5346; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5348 = 6'h24 == _next_rob_state_T_10[5:0] ? rob_uop_36_stale_dst : _GEN_5347; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5349 = 6'h25 == _next_rob_state_T_10[5:0] ? rob_uop_37_stale_dst : _GEN_5348; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5350 = 6'h26 == _next_rob_state_T_10[5:0] ? rob_uop_38_stale_dst : _GEN_5349; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5351 = 6'h27 == _next_rob_state_T_10[5:0] ? rob_uop_39_stale_dst : _GEN_5350; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5352 = 6'h28 == _next_rob_state_T_10[5:0] ? rob_uop_40_stale_dst : _GEN_5351; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5353 = 6'h29 == _next_rob_state_T_10[5:0] ? rob_uop_41_stale_dst : _GEN_5352; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5354 = 6'h2a == _next_rob_state_T_10[5:0] ? rob_uop_42_stale_dst : _GEN_5353; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5355 = 6'h2b == _next_rob_state_T_10[5:0] ? rob_uop_43_stale_dst : _GEN_5354; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5356 = 6'h2c == _next_rob_state_T_10[5:0] ? rob_uop_44_stale_dst : _GEN_5355; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5357 = 6'h2d == _next_rob_state_T_10[5:0] ? rob_uop_45_stale_dst : _GEN_5356; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5358 = 6'h2e == _next_rob_state_T_10[5:0] ? rob_uop_46_stale_dst : _GEN_5357; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5359 = 6'h2f == _next_rob_state_T_10[5:0] ? rob_uop_47_stale_dst : _GEN_5358; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5360 = 6'h30 == _next_rob_state_T_10[5:0] ? rob_uop_48_stale_dst : _GEN_5359; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5361 = 6'h31 == _next_rob_state_T_10[5:0] ? rob_uop_49_stale_dst : _GEN_5360; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5362 = 6'h32 == _next_rob_state_T_10[5:0] ? rob_uop_50_stale_dst : _GEN_5361; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5363 = 6'h33 == _next_rob_state_T_10[5:0] ? rob_uop_51_stale_dst : _GEN_5362; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5364 = 6'h34 == _next_rob_state_T_10[5:0] ? rob_uop_52_stale_dst : _GEN_5363; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5365 = 6'h35 == _next_rob_state_T_10[5:0] ? rob_uop_53_stale_dst : _GEN_5364; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5366 = 6'h36 == _next_rob_state_T_10[5:0] ? rob_uop_54_stale_dst : _GEN_5365; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5367 = 6'h37 == _next_rob_state_T_10[5:0] ? rob_uop_55_stale_dst : _GEN_5366; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5368 = 6'h38 == _next_rob_state_T_10[5:0] ? rob_uop_56_stale_dst : _GEN_5367; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5369 = 6'h39 == _next_rob_state_T_10[5:0] ? rob_uop_57_stale_dst : _GEN_5368; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5370 = 6'h3a == _next_rob_state_T_10[5:0] ? rob_uop_58_stale_dst : _GEN_5369; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5371 = 6'h3b == _next_rob_state_T_10[5:0] ? rob_uop_59_stale_dst : _GEN_5370; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5372 = 6'h3c == _next_rob_state_T_10[5:0] ? rob_uop_60_stale_dst : _GEN_5371; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5373 = 6'h3d == _next_rob_state_T_10[5:0] ? rob_uop_61_stale_dst : _GEN_5372; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_5374 = 6'h3e == _next_rob_state_T_10[5:0] ? rob_uop_62_stale_dst : _GEN_5373; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5377 = 6'h1 == _next_rob_state_T_10[5:0] ? rob_uop_1_arch_dst : rob_uop_0_arch_dst; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5378 = 6'h2 == _next_rob_state_T_10[5:0] ? rob_uop_2_arch_dst : _GEN_5377; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5379 = 6'h3 == _next_rob_state_T_10[5:0] ? rob_uop_3_arch_dst : _GEN_5378; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5380 = 6'h4 == _next_rob_state_T_10[5:0] ? rob_uop_4_arch_dst : _GEN_5379; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5381 = 6'h5 == _next_rob_state_T_10[5:0] ? rob_uop_5_arch_dst : _GEN_5380; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5382 = 6'h6 == _next_rob_state_T_10[5:0] ? rob_uop_6_arch_dst : _GEN_5381; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5383 = 6'h7 == _next_rob_state_T_10[5:0] ? rob_uop_7_arch_dst : _GEN_5382; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5384 = 6'h8 == _next_rob_state_T_10[5:0] ? rob_uop_8_arch_dst : _GEN_5383; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5385 = 6'h9 == _next_rob_state_T_10[5:0] ? rob_uop_9_arch_dst : _GEN_5384; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5386 = 6'ha == _next_rob_state_T_10[5:0] ? rob_uop_10_arch_dst : _GEN_5385; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5387 = 6'hb == _next_rob_state_T_10[5:0] ? rob_uop_11_arch_dst : _GEN_5386; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5388 = 6'hc == _next_rob_state_T_10[5:0] ? rob_uop_12_arch_dst : _GEN_5387; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5389 = 6'hd == _next_rob_state_T_10[5:0] ? rob_uop_13_arch_dst : _GEN_5388; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5390 = 6'he == _next_rob_state_T_10[5:0] ? rob_uop_14_arch_dst : _GEN_5389; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5391 = 6'hf == _next_rob_state_T_10[5:0] ? rob_uop_15_arch_dst : _GEN_5390; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5392 = 6'h10 == _next_rob_state_T_10[5:0] ? rob_uop_16_arch_dst : _GEN_5391; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5393 = 6'h11 == _next_rob_state_T_10[5:0] ? rob_uop_17_arch_dst : _GEN_5392; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5394 = 6'h12 == _next_rob_state_T_10[5:0] ? rob_uop_18_arch_dst : _GEN_5393; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5395 = 6'h13 == _next_rob_state_T_10[5:0] ? rob_uop_19_arch_dst : _GEN_5394; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5396 = 6'h14 == _next_rob_state_T_10[5:0] ? rob_uop_20_arch_dst : _GEN_5395; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5397 = 6'h15 == _next_rob_state_T_10[5:0] ? rob_uop_21_arch_dst : _GEN_5396; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5398 = 6'h16 == _next_rob_state_T_10[5:0] ? rob_uop_22_arch_dst : _GEN_5397; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5399 = 6'h17 == _next_rob_state_T_10[5:0] ? rob_uop_23_arch_dst : _GEN_5398; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5400 = 6'h18 == _next_rob_state_T_10[5:0] ? rob_uop_24_arch_dst : _GEN_5399; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5401 = 6'h19 == _next_rob_state_T_10[5:0] ? rob_uop_25_arch_dst : _GEN_5400; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5402 = 6'h1a == _next_rob_state_T_10[5:0] ? rob_uop_26_arch_dst : _GEN_5401; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5403 = 6'h1b == _next_rob_state_T_10[5:0] ? rob_uop_27_arch_dst : _GEN_5402; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5404 = 6'h1c == _next_rob_state_T_10[5:0] ? rob_uop_28_arch_dst : _GEN_5403; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5405 = 6'h1d == _next_rob_state_T_10[5:0] ? rob_uop_29_arch_dst : _GEN_5404; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5406 = 6'h1e == _next_rob_state_T_10[5:0] ? rob_uop_30_arch_dst : _GEN_5405; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5407 = 6'h1f == _next_rob_state_T_10[5:0] ? rob_uop_31_arch_dst : _GEN_5406; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5408 = 6'h20 == _next_rob_state_T_10[5:0] ? rob_uop_32_arch_dst : _GEN_5407; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5409 = 6'h21 == _next_rob_state_T_10[5:0] ? rob_uop_33_arch_dst : _GEN_5408; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5410 = 6'h22 == _next_rob_state_T_10[5:0] ? rob_uop_34_arch_dst : _GEN_5409; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5411 = 6'h23 == _next_rob_state_T_10[5:0] ? rob_uop_35_arch_dst : _GEN_5410; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5412 = 6'h24 == _next_rob_state_T_10[5:0] ? rob_uop_36_arch_dst : _GEN_5411; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5413 = 6'h25 == _next_rob_state_T_10[5:0] ? rob_uop_37_arch_dst : _GEN_5412; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5414 = 6'h26 == _next_rob_state_T_10[5:0] ? rob_uop_38_arch_dst : _GEN_5413; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5415 = 6'h27 == _next_rob_state_T_10[5:0] ? rob_uop_39_arch_dst : _GEN_5414; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5416 = 6'h28 == _next_rob_state_T_10[5:0] ? rob_uop_40_arch_dst : _GEN_5415; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5417 = 6'h29 == _next_rob_state_T_10[5:0] ? rob_uop_41_arch_dst : _GEN_5416; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5418 = 6'h2a == _next_rob_state_T_10[5:0] ? rob_uop_42_arch_dst : _GEN_5417; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5419 = 6'h2b == _next_rob_state_T_10[5:0] ? rob_uop_43_arch_dst : _GEN_5418; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5420 = 6'h2c == _next_rob_state_T_10[5:0] ? rob_uop_44_arch_dst : _GEN_5419; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5421 = 6'h2d == _next_rob_state_T_10[5:0] ? rob_uop_45_arch_dst : _GEN_5420; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5422 = 6'h2e == _next_rob_state_T_10[5:0] ? rob_uop_46_arch_dst : _GEN_5421; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5423 = 6'h2f == _next_rob_state_T_10[5:0] ? rob_uop_47_arch_dst : _GEN_5422; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5424 = 6'h30 == _next_rob_state_T_10[5:0] ? rob_uop_48_arch_dst : _GEN_5423; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5425 = 6'h31 == _next_rob_state_T_10[5:0] ? rob_uop_49_arch_dst : _GEN_5424; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5426 = 6'h32 == _next_rob_state_T_10[5:0] ? rob_uop_50_arch_dst : _GEN_5425; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5427 = 6'h33 == _next_rob_state_T_10[5:0] ? rob_uop_51_arch_dst : _GEN_5426; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5428 = 6'h34 == _next_rob_state_T_10[5:0] ? rob_uop_52_arch_dst : _GEN_5427; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5429 = 6'h35 == _next_rob_state_T_10[5:0] ? rob_uop_53_arch_dst : _GEN_5428; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5430 = 6'h36 == _next_rob_state_T_10[5:0] ? rob_uop_54_arch_dst : _GEN_5429; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5431 = 6'h37 == _next_rob_state_T_10[5:0] ? rob_uop_55_arch_dst : _GEN_5430; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5432 = 6'h38 == _next_rob_state_T_10[5:0] ? rob_uop_56_arch_dst : _GEN_5431; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5433 = 6'h39 == _next_rob_state_T_10[5:0] ? rob_uop_57_arch_dst : _GEN_5432; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5434 = 6'h3a == _next_rob_state_T_10[5:0] ? rob_uop_58_arch_dst : _GEN_5433; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5435 = 6'h3b == _next_rob_state_T_10[5:0] ? rob_uop_59_arch_dst : _GEN_5434; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5436 = 6'h3c == _next_rob_state_T_10[5:0] ? rob_uop_60_arch_dst : _GEN_5435; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5437 = 6'h3d == _next_rob_state_T_10[5:0] ? rob_uop_61_arch_dst : _GEN_5436; // @[rob.scala 117:{33,33}]
  wire [4:0] _GEN_5438 = 6'h3e == _next_rob_state_T_10[5:0] ? rob_uop_62_arch_dst : _GEN_5437; // @[rob.scala 117:{33,33}]
  wire [6:0] _GEN_7233 = 6'h1 == _next_rob_state_T_13[5:0] ? rob_uop_1_phy_dst : rob_uop_0_phy_dst; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7234 = 6'h2 == _next_rob_state_T_13[5:0] ? rob_uop_2_phy_dst : _GEN_7233; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7235 = 6'h3 == _next_rob_state_T_13[5:0] ? rob_uop_3_phy_dst : _GEN_7234; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7236 = 6'h4 == _next_rob_state_T_13[5:0] ? rob_uop_4_phy_dst : _GEN_7235; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7237 = 6'h5 == _next_rob_state_T_13[5:0] ? rob_uop_5_phy_dst : _GEN_7236; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7238 = 6'h6 == _next_rob_state_T_13[5:0] ? rob_uop_6_phy_dst : _GEN_7237; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7239 = 6'h7 == _next_rob_state_T_13[5:0] ? rob_uop_7_phy_dst : _GEN_7238; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7240 = 6'h8 == _next_rob_state_T_13[5:0] ? rob_uop_8_phy_dst : _GEN_7239; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7241 = 6'h9 == _next_rob_state_T_13[5:0] ? rob_uop_9_phy_dst : _GEN_7240; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7242 = 6'ha == _next_rob_state_T_13[5:0] ? rob_uop_10_phy_dst : _GEN_7241; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7243 = 6'hb == _next_rob_state_T_13[5:0] ? rob_uop_11_phy_dst : _GEN_7242; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7244 = 6'hc == _next_rob_state_T_13[5:0] ? rob_uop_12_phy_dst : _GEN_7243; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7245 = 6'hd == _next_rob_state_T_13[5:0] ? rob_uop_13_phy_dst : _GEN_7244; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7246 = 6'he == _next_rob_state_T_13[5:0] ? rob_uop_14_phy_dst : _GEN_7245; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7247 = 6'hf == _next_rob_state_T_13[5:0] ? rob_uop_15_phy_dst : _GEN_7246; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7248 = 6'h10 == _next_rob_state_T_13[5:0] ? rob_uop_16_phy_dst : _GEN_7247; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7249 = 6'h11 == _next_rob_state_T_13[5:0] ? rob_uop_17_phy_dst : _GEN_7248; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7250 = 6'h12 == _next_rob_state_T_13[5:0] ? rob_uop_18_phy_dst : _GEN_7249; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7251 = 6'h13 == _next_rob_state_T_13[5:0] ? rob_uop_19_phy_dst : _GEN_7250; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7252 = 6'h14 == _next_rob_state_T_13[5:0] ? rob_uop_20_phy_dst : _GEN_7251; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7253 = 6'h15 == _next_rob_state_T_13[5:0] ? rob_uop_21_phy_dst : _GEN_7252; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7254 = 6'h16 == _next_rob_state_T_13[5:0] ? rob_uop_22_phy_dst : _GEN_7253; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7255 = 6'h17 == _next_rob_state_T_13[5:0] ? rob_uop_23_phy_dst : _GEN_7254; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7256 = 6'h18 == _next_rob_state_T_13[5:0] ? rob_uop_24_phy_dst : _GEN_7255; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7257 = 6'h19 == _next_rob_state_T_13[5:0] ? rob_uop_25_phy_dst : _GEN_7256; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7258 = 6'h1a == _next_rob_state_T_13[5:0] ? rob_uop_26_phy_dst : _GEN_7257; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7259 = 6'h1b == _next_rob_state_T_13[5:0] ? rob_uop_27_phy_dst : _GEN_7258; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7260 = 6'h1c == _next_rob_state_T_13[5:0] ? rob_uop_28_phy_dst : _GEN_7259; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7261 = 6'h1d == _next_rob_state_T_13[5:0] ? rob_uop_29_phy_dst : _GEN_7260; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7262 = 6'h1e == _next_rob_state_T_13[5:0] ? rob_uop_30_phy_dst : _GEN_7261; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7263 = 6'h1f == _next_rob_state_T_13[5:0] ? rob_uop_31_phy_dst : _GEN_7262; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7264 = 6'h20 == _next_rob_state_T_13[5:0] ? rob_uop_32_phy_dst : _GEN_7263; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7265 = 6'h21 == _next_rob_state_T_13[5:0] ? rob_uop_33_phy_dst : _GEN_7264; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7266 = 6'h22 == _next_rob_state_T_13[5:0] ? rob_uop_34_phy_dst : _GEN_7265; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7267 = 6'h23 == _next_rob_state_T_13[5:0] ? rob_uop_35_phy_dst : _GEN_7266; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7268 = 6'h24 == _next_rob_state_T_13[5:0] ? rob_uop_36_phy_dst : _GEN_7267; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7269 = 6'h25 == _next_rob_state_T_13[5:0] ? rob_uop_37_phy_dst : _GEN_7268; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7270 = 6'h26 == _next_rob_state_T_13[5:0] ? rob_uop_38_phy_dst : _GEN_7269; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7271 = 6'h27 == _next_rob_state_T_13[5:0] ? rob_uop_39_phy_dst : _GEN_7270; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7272 = 6'h28 == _next_rob_state_T_13[5:0] ? rob_uop_40_phy_dst : _GEN_7271; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7273 = 6'h29 == _next_rob_state_T_13[5:0] ? rob_uop_41_phy_dst : _GEN_7272; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7274 = 6'h2a == _next_rob_state_T_13[5:0] ? rob_uop_42_phy_dst : _GEN_7273; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7275 = 6'h2b == _next_rob_state_T_13[5:0] ? rob_uop_43_phy_dst : _GEN_7274; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7276 = 6'h2c == _next_rob_state_T_13[5:0] ? rob_uop_44_phy_dst : _GEN_7275; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7277 = 6'h2d == _next_rob_state_T_13[5:0] ? rob_uop_45_phy_dst : _GEN_7276; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7278 = 6'h2e == _next_rob_state_T_13[5:0] ? rob_uop_46_phy_dst : _GEN_7277; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7279 = 6'h2f == _next_rob_state_T_13[5:0] ? rob_uop_47_phy_dst : _GEN_7278; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7280 = 6'h30 == _next_rob_state_T_13[5:0] ? rob_uop_48_phy_dst : _GEN_7279; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7281 = 6'h31 == _next_rob_state_T_13[5:0] ? rob_uop_49_phy_dst : _GEN_7280; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7282 = 6'h32 == _next_rob_state_T_13[5:0] ? rob_uop_50_phy_dst : _GEN_7281; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7283 = 6'h33 == _next_rob_state_T_13[5:0] ? rob_uop_51_phy_dst : _GEN_7282; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7284 = 6'h34 == _next_rob_state_T_13[5:0] ? rob_uop_52_phy_dst : _GEN_7283; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7285 = 6'h35 == _next_rob_state_T_13[5:0] ? rob_uop_53_phy_dst : _GEN_7284; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7286 = 6'h36 == _next_rob_state_T_13[5:0] ? rob_uop_54_phy_dst : _GEN_7285; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7287 = 6'h37 == _next_rob_state_T_13[5:0] ? rob_uop_55_phy_dst : _GEN_7286; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7288 = 6'h38 == _next_rob_state_T_13[5:0] ? rob_uop_56_phy_dst : _GEN_7287; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7289 = 6'h39 == _next_rob_state_T_13[5:0] ? rob_uop_57_phy_dst : _GEN_7288; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7290 = 6'h3a == _next_rob_state_T_13[5:0] ? rob_uop_58_phy_dst : _GEN_7289; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7291 = 6'h3b == _next_rob_state_T_13[5:0] ? rob_uop_59_phy_dst : _GEN_7290; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7292 = 6'h3c == _next_rob_state_T_13[5:0] ? rob_uop_60_phy_dst : _GEN_7291; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7293 = 6'h3d == _next_rob_state_T_13[5:0] ? rob_uop_61_phy_dst : _GEN_7292; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7294 = 6'h3e == _next_rob_state_T_13[5:0] ? rob_uop_62_phy_dst : _GEN_7293; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7297 = 6'h1 == _next_rob_state_T_13[5:0] ? rob_uop_1_stale_dst : rob_uop_0_stale_dst; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7298 = 6'h2 == _next_rob_state_T_13[5:0] ? rob_uop_2_stale_dst : _GEN_7297; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7299 = 6'h3 == _next_rob_state_T_13[5:0] ? rob_uop_3_stale_dst : _GEN_7298; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7300 = 6'h4 == _next_rob_state_T_13[5:0] ? rob_uop_4_stale_dst : _GEN_7299; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7301 = 6'h5 == _next_rob_state_T_13[5:0] ? rob_uop_5_stale_dst : _GEN_7300; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7302 = 6'h6 == _next_rob_state_T_13[5:0] ? rob_uop_6_stale_dst : _GEN_7301; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7303 = 6'h7 == _next_rob_state_T_13[5:0] ? rob_uop_7_stale_dst : _GEN_7302; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7304 = 6'h8 == _next_rob_state_T_13[5:0] ? rob_uop_8_stale_dst : _GEN_7303; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7305 = 6'h9 == _next_rob_state_T_13[5:0] ? rob_uop_9_stale_dst : _GEN_7304; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7306 = 6'ha == _next_rob_state_T_13[5:0] ? rob_uop_10_stale_dst : _GEN_7305; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7307 = 6'hb == _next_rob_state_T_13[5:0] ? rob_uop_11_stale_dst : _GEN_7306; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7308 = 6'hc == _next_rob_state_T_13[5:0] ? rob_uop_12_stale_dst : _GEN_7307; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7309 = 6'hd == _next_rob_state_T_13[5:0] ? rob_uop_13_stale_dst : _GEN_7308; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7310 = 6'he == _next_rob_state_T_13[5:0] ? rob_uop_14_stale_dst : _GEN_7309; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7311 = 6'hf == _next_rob_state_T_13[5:0] ? rob_uop_15_stale_dst : _GEN_7310; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7312 = 6'h10 == _next_rob_state_T_13[5:0] ? rob_uop_16_stale_dst : _GEN_7311; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7313 = 6'h11 == _next_rob_state_T_13[5:0] ? rob_uop_17_stale_dst : _GEN_7312; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7314 = 6'h12 == _next_rob_state_T_13[5:0] ? rob_uop_18_stale_dst : _GEN_7313; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7315 = 6'h13 == _next_rob_state_T_13[5:0] ? rob_uop_19_stale_dst : _GEN_7314; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7316 = 6'h14 == _next_rob_state_T_13[5:0] ? rob_uop_20_stale_dst : _GEN_7315; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7317 = 6'h15 == _next_rob_state_T_13[5:0] ? rob_uop_21_stale_dst : _GEN_7316; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7318 = 6'h16 == _next_rob_state_T_13[5:0] ? rob_uop_22_stale_dst : _GEN_7317; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7319 = 6'h17 == _next_rob_state_T_13[5:0] ? rob_uop_23_stale_dst : _GEN_7318; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7320 = 6'h18 == _next_rob_state_T_13[5:0] ? rob_uop_24_stale_dst : _GEN_7319; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7321 = 6'h19 == _next_rob_state_T_13[5:0] ? rob_uop_25_stale_dst : _GEN_7320; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7322 = 6'h1a == _next_rob_state_T_13[5:0] ? rob_uop_26_stale_dst : _GEN_7321; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7323 = 6'h1b == _next_rob_state_T_13[5:0] ? rob_uop_27_stale_dst : _GEN_7322; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7324 = 6'h1c == _next_rob_state_T_13[5:0] ? rob_uop_28_stale_dst : _GEN_7323; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7325 = 6'h1d == _next_rob_state_T_13[5:0] ? rob_uop_29_stale_dst : _GEN_7324; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7326 = 6'h1e == _next_rob_state_T_13[5:0] ? rob_uop_30_stale_dst : _GEN_7325; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7327 = 6'h1f == _next_rob_state_T_13[5:0] ? rob_uop_31_stale_dst : _GEN_7326; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7328 = 6'h20 == _next_rob_state_T_13[5:0] ? rob_uop_32_stale_dst : _GEN_7327; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7329 = 6'h21 == _next_rob_state_T_13[5:0] ? rob_uop_33_stale_dst : _GEN_7328; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7330 = 6'h22 == _next_rob_state_T_13[5:0] ? rob_uop_34_stale_dst : _GEN_7329; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7331 = 6'h23 == _next_rob_state_T_13[5:0] ? rob_uop_35_stale_dst : _GEN_7330; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7332 = 6'h24 == _next_rob_state_T_13[5:0] ? rob_uop_36_stale_dst : _GEN_7331; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7333 = 6'h25 == _next_rob_state_T_13[5:0] ? rob_uop_37_stale_dst : _GEN_7332; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7334 = 6'h26 == _next_rob_state_T_13[5:0] ? rob_uop_38_stale_dst : _GEN_7333; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7335 = 6'h27 == _next_rob_state_T_13[5:0] ? rob_uop_39_stale_dst : _GEN_7334; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7336 = 6'h28 == _next_rob_state_T_13[5:0] ? rob_uop_40_stale_dst : _GEN_7335; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7337 = 6'h29 == _next_rob_state_T_13[5:0] ? rob_uop_41_stale_dst : _GEN_7336; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7338 = 6'h2a == _next_rob_state_T_13[5:0] ? rob_uop_42_stale_dst : _GEN_7337; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7339 = 6'h2b == _next_rob_state_T_13[5:0] ? rob_uop_43_stale_dst : _GEN_7338; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7340 = 6'h2c == _next_rob_state_T_13[5:0] ? rob_uop_44_stale_dst : _GEN_7339; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7341 = 6'h2d == _next_rob_state_T_13[5:0] ? rob_uop_45_stale_dst : _GEN_7340; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7342 = 6'h2e == _next_rob_state_T_13[5:0] ? rob_uop_46_stale_dst : _GEN_7341; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7343 = 6'h2f == _next_rob_state_T_13[5:0] ? rob_uop_47_stale_dst : _GEN_7342; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7344 = 6'h30 == _next_rob_state_T_13[5:0] ? rob_uop_48_stale_dst : _GEN_7343; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7345 = 6'h31 == _next_rob_state_T_13[5:0] ? rob_uop_49_stale_dst : _GEN_7344; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7346 = 6'h32 == _next_rob_state_T_13[5:0] ? rob_uop_50_stale_dst : _GEN_7345; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7347 = 6'h33 == _next_rob_state_T_13[5:0] ? rob_uop_51_stale_dst : _GEN_7346; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7348 = 6'h34 == _next_rob_state_T_13[5:0] ? rob_uop_52_stale_dst : _GEN_7347; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7349 = 6'h35 == _next_rob_state_T_13[5:0] ? rob_uop_53_stale_dst : _GEN_7348; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7350 = 6'h36 == _next_rob_state_T_13[5:0] ? rob_uop_54_stale_dst : _GEN_7349; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7351 = 6'h37 == _next_rob_state_T_13[5:0] ? rob_uop_55_stale_dst : _GEN_7350; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7352 = 6'h38 == _next_rob_state_T_13[5:0] ? rob_uop_56_stale_dst : _GEN_7351; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7353 = 6'h39 == _next_rob_state_T_13[5:0] ? rob_uop_57_stale_dst : _GEN_7352; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7354 = 6'h3a == _next_rob_state_T_13[5:0] ? rob_uop_58_stale_dst : _GEN_7353; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7355 = 6'h3b == _next_rob_state_T_13[5:0] ? rob_uop_59_stale_dst : _GEN_7354; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7356 = 6'h3c == _next_rob_state_T_13[5:0] ? rob_uop_60_stale_dst : _GEN_7355; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7357 = 6'h3d == _next_rob_state_T_13[5:0] ? rob_uop_61_stale_dst : _GEN_7356; // @[rob.scala 118:{33,33}]
  wire [6:0] _GEN_7358 = 6'h3e == _next_rob_state_T_13[5:0] ? rob_uop_62_stale_dst : _GEN_7357; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7361 = 6'h1 == _next_rob_state_T_13[5:0] ? rob_uop_1_arch_dst : rob_uop_0_arch_dst; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7362 = 6'h2 == _next_rob_state_T_13[5:0] ? rob_uop_2_arch_dst : _GEN_7361; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7363 = 6'h3 == _next_rob_state_T_13[5:0] ? rob_uop_3_arch_dst : _GEN_7362; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7364 = 6'h4 == _next_rob_state_T_13[5:0] ? rob_uop_4_arch_dst : _GEN_7363; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7365 = 6'h5 == _next_rob_state_T_13[5:0] ? rob_uop_5_arch_dst : _GEN_7364; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7366 = 6'h6 == _next_rob_state_T_13[5:0] ? rob_uop_6_arch_dst : _GEN_7365; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7367 = 6'h7 == _next_rob_state_T_13[5:0] ? rob_uop_7_arch_dst : _GEN_7366; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7368 = 6'h8 == _next_rob_state_T_13[5:0] ? rob_uop_8_arch_dst : _GEN_7367; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7369 = 6'h9 == _next_rob_state_T_13[5:0] ? rob_uop_9_arch_dst : _GEN_7368; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7370 = 6'ha == _next_rob_state_T_13[5:0] ? rob_uop_10_arch_dst : _GEN_7369; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7371 = 6'hb == _next_rob_state_T_13[5:0] ? rob_uop_11_arch_dst : _GEN_7370; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7372 = 6'hc == _next_rob_state_T_13[5:0] ? rob_uop_12_arch_dst : _GEN_7371; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7373 = 6'hd == _next_rob_state_T_13[5:0] ? rob_uop_13_arch_dst : _GEN_7372; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7374 = 6'he == _next_rob_state_T_13[5:0] ? rob_uop_14_arch_dst : _GEN_7373; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7375 = 6'hf == _next_rob_state_T_13[5:0] ? rob_uop_15_arch_dst : _GEN_7374; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7376 = 6'h10 == _next_rob_state_T_13[5:0] ? rob_uop_16_arch_dst : _GEN_7375; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7377 = 6'h11 == _next_rob_state_T_13[5:0] ? rob_uop_17_arch_dst : _GEN_7376; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7378 = 6'h12 == _next_rob_state_T_13[5:0] ? rob_uop_18_arch_dst : _GEN_7377; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7379 = 6'h13 == _next_rob_state_T_13[5:0] ? rob_uop_19_arch_dst : _GEN_7378; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7380 = 6'h14 == _next_rob_state_T_13[5:0] ? rob_uop_20_arch_dst : _GEN_7379; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7381 = 6'h15 == _next_rob_state_T_13[5:0] ? rob_uop_21_arch_dst : _GEN_7380; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7382 = 6'h16 == _next_rob_state_T_13[5:0] ? rob_uop_22_arch_dst : _GEN_7381; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7383 = 6'h17 == _next_rob_state_T_13[5:0] ? rob_uop_23_arch_dst : _GEN_7382; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7384 = 6'h18 == _next_rob_state_T_13[5:0] ? rob_uop_24_arch_dst : _GEN_7383; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7385 = 6'h19 == _next_rob_state_T_13[5:0] ? rob_uop_25_arch_dst : _GEN_7384; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7386 = 6'h1a == _next_rob_state_T_13[5:0] ? rob_uop_26_arch_dst : _GEN_7385; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7387 = 6'h1b == _next_rob_state_T_13[5:0] ? rob_uop_27_arch_dst : _GEN_7386; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7388 = 6'h1c == _next_rob_state_T_13[5:0] ? rob_uop_28_arch_dst : _GEN_7387; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7389 = 6'h1d == _next_rob_state_T_13[5:0] ? rob_uop_29_arch_dst : _GEN_7388; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7390 = 6'h1e == _next_rob_state_T_13[5:0] ? rob_uop_30_arch_dst : _GEN_7389; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7391 = 6'h1f == _next_rob_state_T_13[5:0] ? rob_uop_31_arch_dst : _GEN_7390; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7392 = 6'h20 == _next_rob_state_T_13[5:0] ? rob_uop_32_arch_dst : _GEN_7391; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7393 = 6'h21 == _next_rob_state_T_13[5:0] ? rob_uop_33_arch_dst : _GEN_7392; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7394 = 6'h22 == _next_rob_state_T_13[5:0] ? rob_uop_34_arch_dst : _GEN_7393; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7395 = 6'h23 == _next_rob_state_T_13[5:0] ? rob_uop_35_arch_dst : _GEN_7394; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7396 = 6'h24 == _next_rob_state_T_13[5:0] ? rob_uop_36_arch_dst : _GEN_7395; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7397 = 6'h25 == _next_rob_state_T_13[5:0] ? rob_uop_37_arch_dst : _GEN_7396; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7398 = 6'h26 == _next_rob_state_T_13[5:0] ? rob_uop_38_arch_dst : _GEN_7397; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7399 = 6'h27 == _next_rob_state_T_13[5:0] ? rob_uop_39_arch_dst : _GEN_7398; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7400 = 6'h28 == _next_rob_state_T_13[5:0] ? rob_uop_40_arch_dst : _GEN_7399; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7401 = 6'h29 == _next_rob_state_T_13[5:0] ? rob_uop_41_arch_dst : _GEN_7400; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7402 = 6'h2a == _next_rob_state_T_13[5:0] ? rob_uop_42_arch_dst : _GEN_7401; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7403 = 6'h2b == _next_rob_state_T_13[5:0] ? rob_uop_43_arch_dst : _GEN_7402; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7404 = 6'h2c == _next_rob_state_T_13[5:0] ? rob_uop_44_arch_dst : _GEN_7403; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7405 = 6'h2d == _next_rob_state_T_13[5:0] ? rob_uop_45_arch_dst : _GEN_7404; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7406 = 6'h2e == _next_rob_state_T_13[5:0] ? rob_uop_46_arch_dst : _GEN_7405; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7407 = 6'h2f == _next_rob_state_T_13[5:0] ? rob_uop_47_arch_dst : _GEN_7406; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7408 = 6'h30 == _next_rob_state_T_13[5:0] ? rob_uop_48_arch_dst : _GEN_7407; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7409 = 6'h31 == _next_rob_state_T_13[5:0] ? rob_uop_49_arch_dst : _GEN_7408; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7410 = 6'h32 == _next_rob_state_T_13[5:0] ? rob_uop_50_arch_dst : _GEN_7409; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7411 = 6'h33 == _next_rob_state_T_13[5:0] ? rob_uop_51_arch_dst : _GEN_7410; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7412 = 6'h34 == _next_rob_state_T_13[5:0] ? rob_uop_52_arch_dst : _GEN_7411; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7413 = 6'h35 == _next_rob_state_T_13[5:0] ? rob_uop_53_arch_dst : _GEN_7412; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7414 = 6'h36 == _next_rob_state_T_13[5:0] ? rob_uop_54_arch_dst : _GEN_7413; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7415 = 6'h37 == _next_rob_state_T_13[5:0] ? rob_uop_55_arch_dst : _GEN_7414; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7416 = 6'h38 == _next_rob_state_T_13[5:0] ? rob_uop_56_arch_dst : _GEN_7415; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7417 = 6'h39 == _next_rob_state_T_13[5:0] ? rob_uop_57_arch_dst : _GEN_7416; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7418 = 6'h3a == _next_rob_state_T_13[5:0] ? rob_uop_58_arch_dst : _GEN_7417; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7419 = 6'h3b == _next_rob_state_T_13[5:0] ? rob_uop_59_arch_dst : _GEN_7418; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7420 = 6'h3c == _next_rob_state_T_13[5:0] ? rob_uop_60_arch_dst : _GEN_7419; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7421 = 6'h3d == _next_rob_state_T_13[5:0] ? rob_uop_61_arch_dst : _GEN_7420; // @[rob.scala 118:{33,33}]
  wire [4:0] _GEN_7422 = 6'h3e == _next_rob_state_T_13[5:0] ? rob_uop_62_arch_dst : _GEN_7421; // @[rob.scala 118:{33,33}]
  wire [31:0] _GEN_8704 = 6'h0 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_0_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8705 = 6'h1 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_1_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8706 = 6'h2 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_2_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8707 = 6'h3 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_3_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8708 = 6'h4 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_4_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8709 = 6'h5 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_5_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8710 = 6'h6 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_6_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8711 = 6'h7 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_7_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8712 = 6'h8 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_8_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8713 = 6'h9 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_9_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8714 = 6'ha == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_10_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8715 = 6'hb == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_11_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8716 = 6'hc == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_12_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8717 = 6'hd == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_13_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8718 = 6'he == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_14_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8719 = 6'hf == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_15_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8720 = 6'h10 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_16_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8721 = 6'h11 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_17_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8722 = 6'h12 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_18_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8723 = 6'h13 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_19_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8724 = 6'h14 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_20_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8725 = 6'h15 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_21_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8726 = 6'h16 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_22_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8727 = 6'h17 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_23_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8728 = 6'h18 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_24_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8729 = 6'h19 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_25_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8730 = 6'h1a == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_26_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8731 = 6'h1b == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_27_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8732 = 6'h1c == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_28_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8733 = 6'h1d == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_29_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8734 = 6'h1e == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_30_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8735 = 6'h1f == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_31_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8736 = 6'h20 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_32_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8737 = 6'h21 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_33_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8738 = 6'h22 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_34_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8739 = 6'h23 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_35_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8740 = 6'h24 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_36_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8741 = 6'h25 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_37_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8742 = 6'h26 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_38_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8743 = 6'h27 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_39_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8744 = 6'h28 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_40_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8745 = 6'h29 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_41_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8746 = 6'h2a == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_42_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8747 = 6'h2b == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_43_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8748 = 6'h2c == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_44_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8749 = 6'h2d == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_45_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8750 = 6'h2e == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_46_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8751 = 6'h2f == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_47_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8752 = 6'h30 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_48_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8753 = 6'h31 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_49_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8754 = 6'h32 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_50_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8755 = 6'h33 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_51_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8756 = 6'h34 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_52_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8757 = 6'h35 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_53_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8758 = 6'h36 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_54_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8759 = 6'h37 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_55_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8760 = 6'h38 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_56_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8761 = 6'h39 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_57_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8762 = 6'h3a == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_58_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8763 = 6'h3b == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_59_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8764 = 6'h3c == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_60_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8765 = 6'h3d == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_61_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8766 = 6'h3e == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_62_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8767 = 6'h3f == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_pc : rob_uop_63_pc; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8768 = 6'h0 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_0_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8769 = 6'h1 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_1_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8770 = 6'h2 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_2_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8771 = 6'h3 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_3_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8772 = 6'h4 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_4_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8773 = 6'h5 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_5_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8774 = 6'h6 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_6_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8775 = 6'h7 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_7_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8776 = 6'h8 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_8_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8777 = 6'h9 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_9_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8778 = 6'ha == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_10_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8779 = 6'hb == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_11_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8780 = 6'hc == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_12_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8781 = 6'hd == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_13_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8782 = 6'he == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_14_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8783 = 6'hf == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_15_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8784 = 6'h10 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_16_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8785 = 6'h11 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_17_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8786 = 6'h12 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_18_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8787 = 6'h13 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_19_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8788 = 6'h14 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_20_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8789 = 6'h15 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_21_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8790 = 6'h16 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_22_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8791 = 6'h17 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_23_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8792 = 6'h18 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_24_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8793 = 6'h19 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_25_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8794 = 6'h1a == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_26_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8795 = 6'h1b == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_27_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8796 = 6'h1c == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_28_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8797 = 6'h1d == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_29_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8798 = 6'h1e == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_30_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8799 = 6'h1f == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_31_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8800 = 6'h20 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_32_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8801 = 6'h21 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_33_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8802 = 6'h22 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_34_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8803 = 6'h23 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_35_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8804 = 6'h24 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_36_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8805 = 6'h25 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_37_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8806 = 6'h26 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_38_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8807 = 6'h27 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_39_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8808 = 6'h28 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_40_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8809 = 6'h29 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_41_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8810 = 6'h2a == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_42_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8811 = 6'h2b == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_43_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8812 = 6'h2c == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_44_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8813 = 6'h2d == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_45_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8814 = 6'h2e == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_46_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8815 = 6'h2f == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_47_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8816 = 6'h30 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_48_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8817 = 6'h31 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_49_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8818 = 6'h32 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_50_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8819 = 6'h33 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_51_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8820 = 6'h34 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_52_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8821 = 6'h35 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_53_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8822 = 6'h36 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_54_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8823 = 6'h37 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_55_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8824 = 6'h38 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_56_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8825 = 6'h39 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_57_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8826 = 6'h3a == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_58_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8827 = 6'h3b == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_59_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8828 = 6'h3c == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_60_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8829 = 6'h3d == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_61_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8830 = 6'h3e == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_62_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [31:0] _GEN_8831 = 6'h3f == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_inst : rob_uop_63_inst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8832 = 6'h0 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_0_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8833 = 6'h1 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_1_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8834 = 6'h2 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_2_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8835 = 6'h3 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_3_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8836 = 6'h4 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_4_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8837 = 6'h5 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_5_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8838 = 6'h6 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_6_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8839 = 6'h7 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_7_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8840 = 6'h8 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_8_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8841 = 6'h9 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_9_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8842 = 6'ha == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_10_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8843 = 6'hb == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_11_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8844 = 6'hc == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_12_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8845 = 6'hd == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_13_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8846 = 6'he == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_14_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8847 = 6'hf == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_15_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8848 = 6'h10 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_16_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8849 = 6'h11 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_17_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8850 = 6'h12 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_18_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8851 = 6'h13 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_19_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8852 = 6'h14 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_20_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8853 = 6'h15 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_21_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8854 = 6'h16 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_22_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8855 = 6'h17 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_23_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8856 = 6'h18 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_24_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8857 = 6'h19 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_25_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8858 = 6'h1a == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_26_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8859 = 6'h1b == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_27_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8860 = 6'h1c == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_28_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8861 = 6'h1d == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_29_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8862 = 6'h1e == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_30_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8863 = 6'h1f == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_31_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8864 = 6'h20 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_32_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8865 = 6'h21 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_33_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8866 = 6'h22 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_34_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8867 = 6'h23 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_35_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8868 = 6'h24 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_36_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8869 = 6'h25 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_37_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8870 = 6'h26 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_38_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8871 = 6'h27 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_39_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8872 = 6'h28 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_40_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8873 = 6'h29 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_41_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8874 = 6'h2a == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_42_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8875 = 6'h2b == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_43_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8876 = 6'h2c == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_44_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8877 = 6'h2d == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_45_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8878 = 6'h2e == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_46_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8879 = 6'h2f == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_47_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8880 = 6'h30 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_48_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8881 = 6'h31 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_49_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8882 = 6'h32 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_50_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8883 = 6'h33 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_51_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8884 = 6'h34 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_52_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8885 = 6'h35 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_53_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8886 = 6'h36 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_54_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8887 = 6'h37 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_55_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8888 = 6'h38 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_56_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8889 = 6'h39 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_57_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8890 = 6'h3a == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_58_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8891 = 6'h3b == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_59_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8892 = 6'h3c == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_60_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8893 = 6'h3d == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_61_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8894 = 6'h3e == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_62_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_8895 = 6'h3f == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_func_code : rob_uop_63_func_code; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9216 = 6'h0 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_0_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9217 = 6'h1 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_1_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9218 = 6'h2 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_2_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9219 = 6'h3 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_3_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9220 = 6'h4 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_4_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9221 = 6'h5 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_5_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9222 = 6'h6 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_6_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9223 = 6'h7 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_7_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9224 = 6'h8 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_8_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9225 = 6'h9 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_9_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9226 = 6'ha == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_10_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9227 = 6'hb == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_11_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9228 = 6'hc == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_12_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9229 = 6'hd == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_13_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9230 = 6'he == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_14_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9231 = 6'hf == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_15_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9232 = 6'h10 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_16_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9233 = 6'h11 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_17_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9234 = 6'h12 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_18_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9235 = 6'h13 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_19_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9236 = 6'h14 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_20_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9237 = 6'h15 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_21_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9238 = 6'h16 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_22_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9239 = 6'h17 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_23_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9240 = 6'h18 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_24_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9241 = 6'h19 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_25_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9242 = 6'h1a == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_26_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9243 = 6'h1b == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_27_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9244 = 6'h1c == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_28_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9245 = 6'h1d == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_29_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9246 = 6'h1e == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_30_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9247 = 6'h1f == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_31_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9248 = 6'h20 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_32_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9249 = 6'h21 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_33_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9250 = 6'h22 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_34_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9251 = 6'h23 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_35_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9252 = 6'h24 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_36_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9253 = 6'h25 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_37_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9254 = 6'h26 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_38_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9255 = 6'h27 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_39_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9256 = 6'h28 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_40_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9257 = 6'h29 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_41_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9258 = 6'h2a == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_42_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9259 = 6'h2b == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_43_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9260 = 6'h2c == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_44_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9261 = 6'h2d == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_45_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9262 = 6'h2e == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_46_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9263 = 6'h2f == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_47_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9264 = 6'h30 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_48_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9265 = 6'h31 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_49_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9266 = 6'h32 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_50_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9267 = 6'h33 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_51_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9268 = 6'h34 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_52_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9269 = 6'h35 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_53_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9270 = 6'h36 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_54_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9271 = 6'h37 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_55_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9272 = 6'h38 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_56_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9273 = 6'h39 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_57_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9274 = 6'h3a == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_58_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9275 = 6'h3b == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_59_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9276 = 6'h3c == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_60_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9277 = 6'h3d == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_61_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9278 = 6'h3e == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_62_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9279 = 6'h3f == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_phy_dst : rob_uop_63_phy_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9280 = 6'h0 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_0_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9281 = 6'h1 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_1_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9282 = 6'h2 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_2_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9283 = 6'h3 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_3_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9284 = 6'h4 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_4_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9285 = 6'h5 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_5_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9286 = 6'h6 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_6_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9287 = 6'h7 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_7_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9288 = 6'h8 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_8_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9289 = 6'h9 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_9_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9290 = 6'ha == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_10_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9291 = 6'hb == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_11_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9292 = 6'hc == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_12_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9293 = 6'hd == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_13_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9294 = 6'he == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_14_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9295 = 6'hf == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_15_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9296 = 6'h10 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_16_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9297 = 6'h11 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_17_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9298 = 6'h12 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_18_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9299 = 6'h13 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_19_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9300 = 6'h14 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_20_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9301 = 6'h15 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_21_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9302 = 6'h16 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_22_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9303 = 6'h17 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_23_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9304 = 6'h18 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_24_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9305 = 6'h19 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_25_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9306 = 6'h1a == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_26_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9307 = 6'h1b == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_27_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9308 = 6'h1c == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_28_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9309 = 6'h1d == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_29_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9310 = 6'h1e == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_30_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9311 = 6'h1f == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_31_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9312 = 6'h20 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_32_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9313 = 6'h21 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_33_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9314 = 6'h22 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_34_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9315 = 6'h23 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_35_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9316 = 6'h24 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_36_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9317 = 6'h25 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_37_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9318 = 6'h26 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_38_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9319 = 6'h27 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_39_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9320 = 6'h28 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_40_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9321 = 6'h29 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_41_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9322 = 6'h2a == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_42_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9323 = 6'h2b == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_43_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9324 = 6'h2c == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_44_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9325 = 6'h2d == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_45_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9326 = 6'h2e == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_46_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9327 = 6'h2f == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_47_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9328 = 6'h30 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_48_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9329 = 6'h31 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_49_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9330 = 6'h32 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_50_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9331 = 6'h33 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_51_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9332 = 6'h34 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_52_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9333 = 6'h35 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_53_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9334 = 6'h36 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_54_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9335 = 6'h37 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_55_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9336 = 6'h38 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_56_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9337 = 6'h39 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_57_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9338 = 6'h3a == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_58_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9339 = 6'h3b == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_59_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9340 = 6'h3c == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_60_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9341 = 6'h3d == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_61_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9342 = 6'h3e == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_62_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [6:0] _GEN_9343 = 6'h3f == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_stale_dst : rob_uop_63_stale_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9344 = 6'h0 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_0_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9345 = 6'h1 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_1_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9346 = 6'h2 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_2_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9347 = 6'h3 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_3_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9348 = 6'h4 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_4_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9349 = 6'h5 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_5_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9350 = 6'h6 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_6_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9351 = 6'h7 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_7_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9352 = 6'h8 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_8_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9353 = 6'h9 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_9_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9354 = 6'ha == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_10_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9355 = 6'hb == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_11_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9356 = 6'hc == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_12_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9357 = 6'hd == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_13_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9358 = 6'he == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_14_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9359 = 6'hf == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_15_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9360 = 6'h10 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_16_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9361 = 6'h11 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_17_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9362 = 6'h12 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_18_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9363 = 6'h13 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_19_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9364 = 6'h14 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_20_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9365 = 6'h15 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_21_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9366 = 6'h16 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_22_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9367 = 6'h17 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_23_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9368 = 6'h18 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_24_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9369 = 6'h19 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_25_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9370 = 6'h1a == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_26_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9371 = 6'h1b == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_27_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9372 = 6'h1c == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_28_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9373 = 6'h1d == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_29_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9374 = 6'h1e == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_30_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9375 = 6'h1f == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_31_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9376 = 6'h20 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_32_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9377 = 6'h21 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_33_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9378 = 6'h22 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_34_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9379 = 6'h23 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_35_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9380 = 6'h24 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_36_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9381 = 6'h25 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_37_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9382 = 6'h26 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_38_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9383 = 6'h27 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_39_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9384 = 6'h28 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_40_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9385 = 6'h29 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_41_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9386 = 6'h2a == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_42_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9387 = 6'h2b == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_43_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9388 = 6'h2c == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_44_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9389 = 6'h2d == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_45_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9390 = 6'h2e == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_46_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9391 = 6'h2f == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_47_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9392 = 6'h30 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_48_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9393 = 6'h31 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_49_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9394 = 6'h32 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_50_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9395 = 6'h33 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_51_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9396 = 6'h34 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_52_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9397 = 6'h35 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_53_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9398 = 6'h36 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_54_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9399 = 6'h37 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_55_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9400 = 6'h38 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_56_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9401 = 6'h39 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_57_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9402 = 6'h3a == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_58_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9403 = 6'h3b == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_59_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9404 = 6'h3c == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_60_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9405 = 6'h3d == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_61_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9406 = 6'h3e == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_62_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_9407 = 6'h3f == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_arch_dst : rob_uop_63_arch_dst; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10048 = 6'h0 == allocate_ptr[5:0] ? 64'h0 : rob_uop_0_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10049 = 6'h1 == allocate_ptr[5:0] ? 64'h0 : rob_uop_1_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10050 = 6'h2 == allocate_ptr[5:0] ? 64'h0 : rob_uop_2_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10051 = 6'h3 == allocate_ptr[5:0] ? 64'h0 : rob_uop_3_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10052 = 6'h4 == allocate_ptr[5:0] ? 64'h0 : rob_uop_4_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10053 = 6'h5 == allocate_ptr[5:0] ? 64'h0 : rob_uop_5_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10054 = 6'h6 == allocate_ptr[5:0] ? 64'h0 : rob_uop_6_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10055 = 6'h7 == allocate_ptr[5:0] ? 64'h0 : rob_uop_7_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10056 = 6'h8 == allocate_ptr[5:0] ? 64'h0 : rob_uop_8_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10057 = 6'h9 == allocate_ptr[5:0] ? 64'h0 : rob_uop_9_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10058 = 6'ha == allocate_ptr[5:0] ? 64'h0 : rob_uop_10_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10059 = 6'hb == allocate_ptr[5:0] ? 64'h0 : rob_uop_11_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10060 = 6'hc == allocate_ptr[5:0] ? 64'h0 : rob_uop_12_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10061 = 6'hd == allocate_ptr[5:0] ? 64'h0 : rob_uop_13_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10062 = 6'he == allocate_ptr[5:0] ? 64'h0 : rob_uop_14_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10063 = 6'hf == allocate_ptr[5:0] ? 64'h0 : rob_uop_15_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10064 = 6'h10 == allocate_ptr[5:0] ? 64'h0 : rob_uop_16_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10065 = 6'h11 == allocate_ptr[5:0] ? 64'h0 : rob_uop_17_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10066 = 6'h12 == allocate_ptr[5:0] ? 64'h0 : rob_uop_18_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10067 = 6'h13 == allocate_ptr[5:0] ? 64'h0 : rob_uop_19_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10068 = 6'h14 == allocate_ptr[5:0] ? 64'h0 : rob_uop_20_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10069 = 6'h15 == allocate_ptr[5:0] ? 64'h0 : rob_uop_21_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10070 = 6'h16 == allocate_ptr[5:0] ? 64'h0 : rob_uop_22_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10071 = 6'h17 == allocate_ptr[5:0] ? 64'h0 : rob_uop_23_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10072 = 6'h18 == allocate_ptr[5:0] ? 64'h0 : rob_uop_24_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10073 = 6'h19 == allocate_ptr[5:0] ? 64'h0 : rob_uop_25_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10074 = 6'h1a == allocate_ptr[5:0] ? 64'h0 : rob_uop_26_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10075 = 6'h1b == allocate_ptr[5:0] ? 64'h0 : rob_uop_27_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10076 = 6'h1c == allocate_ptr[5:0] ? 64'h0 : rob_uop_28_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10077 = 6'h1d == allocate_ptr[5:0] ? 64'h0 : rob_uop_29_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10078 = 6'h1e == allocate_ptr[5:0] ? 64'h0 : rob_uop_30_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10079 = 6'h1f == allocate_ptr[5:0] ? 64'h0 : rob_uop_31_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10080 = 6'h20 == allocate_ptr[5:0] ? 64'h0 : rob_uop_32_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10081 = 6'h21 == allocate_ptr[5:0] ? 64'h0 : rob_uop_33_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10082 = 6'h22 == allocate_ptr[5:0] ? 64'h0 : rob_uop_34_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10083 = 6'h23 == allocate_ptr[5:0] ? 64'h0 : rob_uop_35_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10084 = 6'h24 == allocate_ptr[5:0] ? 64'h0 : rob_uop_36_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10085 = 6'h25 == allocate_ptr[5:0] ? 64'h0 : rob_uop_37_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10086 = 6'h26 == allocate_ptr[5:0] ? 64'h0 : rob_uop_38_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10087 = 6'h27 == allocate_ptr[5:0] ? 64'h0 : rob_uop_39_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10088 = 6'h28 == allocate_ptr[5:0] ? 64'h0 : rob_uop_40_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10089 = 6'h29 == allocate_ptr[5:0] ? 64'h0 : rob_uop_41_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10090 = 6'h2a == allocate_ptr[5:0] ? 64'h0 : rob_uop_42_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10091 = 6'h2b == allocate_ptr[5:0] ? 64'h0 : rob_uop_43_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10092 = 6'h2c == allocate_ptr[5:0] ? 64'h0 : rob_uop_44_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10093 = 6'h2d == allocate_ptr[5:0] ? 64'h0 : rob_uop_45_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10094 = 6'h2e == allocate_ptr[5:0] ? 64'h0 : rob_uop_46_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10095 = 6'h2f == allocate_ptr[5:0] ? 64'h0 : rob_uop_47_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10096 = 6'h30 == allocate_ptr[5:0] ? 64'h0 : rob_uop_48_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10097 = 6'h31 == allocate_ptr[5:0] ? 64'h0 : rob_uop_49_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10098 = 6'h32 == allocate_ptr[5:0] ? 64'h0 : rob_uop_50_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10099 = 6'h33 == allocate_ptr[5:0] ? 64'h0 : rob_uop_51_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10100 = 6'h34 == allocate_ptr[5:0] ? 64'h0 : rob_uop_52_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10101 = 6'h35 == allocate_ptr[5:0] ? 64'h0 : rob_uop_53_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10102 = 6'h36 == allocate_ptr[5:0] ? 64'h0 : rob_uop_54_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10103 = 6'h37 == allocate_ptr[5:0] ? 64'h0 : rob_uop_55_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10104 = 6'h38 == allocate_ptr[5:0] ? 64'h0 : rob_uop_56_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10105 = 6'h39 == allocate_ptr[5:0] ? 64'h0 : rob_uop_57_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10106 = 6'h3a == allocate_ptr[5:0] ? 64'h0 : rob_uop_58_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10107 = 6'h3b == allocate_ptr[5:0] ? 64'h0 : rob_uop_59_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10108 = 6'h3c == allocate_ptr[5:0] ? 64'h0 : rob_uop_60_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10109 = 6'h3d == allocate_ptr[5:0] ? 64'h0 : rob_uop_61_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10110 = 6'h3e == allocate_ptr[5:0] ? 64'h0 : rob_uop_62_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10111 = 6'h3f == allocate_ptr[5:0] ? 64'h0 : rob_uop_63_dst_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10112 = 6'h0 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value : rob_uop_0_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10113 = 6'h1 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value : rob_uop_1_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10114 = 6'h2 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value : rob_uop_2_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10115 = 6'h3 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value : rob_uop_3_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10116 = 6'h4 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value : rob_uop_4_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10117 = 6'h5 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value : rob_uop_5_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10118 = 6'h6 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value : rob_uop_6_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10119 = 6'h7 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value : rob_uop_7_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10120 = 6'h8 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value : rob_uop_8_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10121 = 6'h9 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value : rob_uop_9_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10122 = 6'ha == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value : rob_uop_10_src1_value
    ; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10123 = 6'hb == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value : rob_uop_11_src1_value
    ; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10124 = 6'hc == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value : rob_uop_12_src1_value
    ; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10125 = 6'hd == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value : rob_uop_13_src1_value
    ; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10126 = 6'he == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value : rob_uop_14_src1_value
    ; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10127 = 6'hf == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value : rob_uop_15_src1_value
    ; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10128 = 6'h10 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_16_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10129 = 6'h11 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_17_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10130 = 6'h12 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_18_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10131 = 6'h13 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_19_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10132 = 6'h14 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_20_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10133 = 6'h15 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_21_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10134 = 6'h16 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_22_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10135 = 6'h17 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_23_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10136 = 6'h18 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_24_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10137 = 6'h19 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_25_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10138 = 6'h1a == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_26_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10139 = 6'h1b == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_27_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10140 = 6'h1c == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_28_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10141 = 6'h1d == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_29_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10142 = 6'h1e == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_30_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10143 = 6'h1f == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_31_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10144 = 6'h20 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_32_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10145 = 6'h21 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_33_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10146 = 6'h22 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_34_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10147 = 6'h23 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_35_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10148 = 6'h24 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_36_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10149 = 6'h25 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_37_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10150 = 6'h26 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_38_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10151 = 6'h27 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_39_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10152 = 6'h28 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_40_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10153 = 6'h29 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_41_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10154 = 6'h2a == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_42_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10155 = 6'h2b == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_43_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10156 = 6'h2c == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_44_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10157 = 6'h2d == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_45_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10158 = 6'h2e == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_46_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10159 = 6'h2f == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_47_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10160 = 6'h30 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_48_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10161 = 6'h31 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_49_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10162 = 6'h32 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_50_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10163 = 6'h33 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_51_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10164 = 6'h34 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_52_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10165 = 6'h35 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_53_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10166 = 6'h36 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_54_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10167 = 6'h37 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_55_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10168 = 6'h38 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_56_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10169 = 6'h39 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_57_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10170 = 6'h3a == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_58_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10171 = 6'h3b == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_59_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10172 = 6'h3c == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_60_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10173 = 6'h3d == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_61_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10174 = 6'h3e == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_62_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [63:0] _GEN_10175 = 6'h3f == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_src1_value :
    rob_uop_63_src1_value; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10432 = 6'h0 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_0_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10433 = 6'h1 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_1_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10434 = 6'h2 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_2_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10435 = 6'h3 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_3_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10436 = 6'h4 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_4_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10437 = 6'h5 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_5_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10438 = 6'h6 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_6_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10439 = 6'h7 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_7_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10440 = 6'h8 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_8_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10441 = 6'h9 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_9_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10442 = 6'ha == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_10_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10443 = 6'hb == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_11_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10444 = 6'hc == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_12_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10445 = 6'hd == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_13_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10446 = 6'he == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_14_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10447 = 6'hf == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_15_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10448 = 6'h10 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_16_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10449 = 6'h11 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_17_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10450 = 6'h12 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_18_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10451 = 6'h13 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_19_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10452 = 6'h14 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_20_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10453 = 6'h15 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_21_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10454 = 6'h16 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_22_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10455 = 6'h17 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_23_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10456 = 6'h18 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_24_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10457 = 6'h19 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_25_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10458 = 6'h1a == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_26_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10459 = 6'h1b == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_27_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10460 = 6'h1c == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_28_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10461 = 6'h1d == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_29_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10462 = 6'h1e == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_30_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10463 = 6'h1f == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_31_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10464 = 6'h20 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_32_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10465 = 6'h21 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_33_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10466 = 6'h22 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_34_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10467 = 6'h23 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_35_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10468 = 6'h24 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_36_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10469 = 6'h25 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_37_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10470 = 6'h26 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_38_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10471 = 6'h27 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_39_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10472 = 6'h28 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_40_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10473 = 6'h29 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_41_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10474 = 6'h2a == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_42_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10475 = 6'h2b == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_43_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10476 = 6'h2c == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_44_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10477 = 6'h2d == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_45_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10478 = 6'h2e == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_46_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10479 = 6'h2f == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_47_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10480 = 6'h30 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_48_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10481 = 6'h31 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_49_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10482 = 6'h32 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_50_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10483 = 6'h33 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_51_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10484 = 6'h34 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_52_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10485 = 6'h35 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_53_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10486 = 6'h36 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_54_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10487 = 6'h37 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_55_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10488 = 6'h38 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_56_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10489 = 6'h39 == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_57_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10490 = 6'h3a == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_58_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10491 = 6'h3b == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_59_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10492 = 6'h3c == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_60_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10493 = 6'h3d == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_61_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10494 = 6'h3e == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_62_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire [4:0] _GEN_10495 = 6'h3f == allocate_ptr[5:0] ? io_i_rob_allocation_reqs_0_uop_alu_sel : rob_uop_63_alu_sel; // @[rob.scala 126:{31,31} 82:26]
  wire  _GEN_10624 = 6'h0 == allocate_ptr[5:0] | rob_valid_0; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10625 = 6'h1 == allocate_ptr[5:0] | rob_valid_1; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10626 = 6'h2 == allocate_ptr[5:0] | rob_valid_2; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10627 = 6'h3 == allocate_ptr[5:0] | rob_valid_3; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10628 = 6'h4 == allocate_ptr[5:0] | rob_valid_4; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10629 = 6'h5 == allocate_ptr[5:0] | rob_valid_5; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10630 = 6'h6 == allocate_ptr[5:0] | rob_valid_6; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10631 = 6'h7 == allocate_ptr[5:0] | rob_valid_7; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10632 = 6'h8 == allocate_ptr[5:0] | rob_valid_8; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10633 = 6'h9 == allocate_ptr[5:0] | rob_valid_9; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10634 = 6'ha == allocate_ptr[5:0] | rob_valid_10; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10635 = 6'hb == allocate_ptr[5:0] | rob_valid_11; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10636 = 6'hc == allocate_ptr[5:0] | rob_valid_12; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10637 = 6'hd == allocate_ptr[5:0] | rob_valid_13; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10638 = 6'he == allocate_ptr[5:0] | rob_valid_14; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10639 = 6'hf == allocate_ptr[5:0] | rob_valid_15; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10640 = 6'h10 == allocate_ptr[5:0] | rob_valid_16; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10641 = 6'h11 == allocate_ptr[5:0] | rob_valid_17; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10642 = 6'h12 == allocate_ptr[5:0] | rob_valid_18; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10643 = 6'h13 == allocate_ptr[5:0] | rob_valid_19; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10644 = 6'h14 == allocate_ptr[5:0] | rob_valid_20; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10645 = 6'h15 == allocate_ptr[5:0] | rob_valid_21; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10646 = 6'h16 == allocate_ptr[5:0] | rob_valid_22; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10647 = 6'h17 == allocate_ptr[5:0] | rob_valid_23; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10648 = 6'h18 == allocate_ptr[5:0] | rob_valid_24; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10649 = 6'h19 == allocate_ptr[5:0] | rob_valid_25; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10650 = 6'h1a == allocate_ptr[5:0] | rob_valid_26; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10651 = 6'h1b == allocate_ptr[5:0] | rob_valid_27; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10652 = 6'h1c == allocate_ptr[5:0] | rob_valid_28; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10653 = 6'h1d == allocate_ptr[5:0] | rob_valid_29; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10654 = 6'h1e == allocate_ptr[5:0] | rob_valid_30; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10655 = 6'h1f == allocate_ptr[5:0] | rob_valid_31; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10656 = 6'h20 == allocate_ptr[5:0] | rob_valid_32; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10657 = 6'h21 == allocate_ptr[5:0] | rob_valid_33; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10658 = 6'h22 == allocate_ptr[5:0] | rob_valid_34; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10659 = 6'h23 == allocate_ptr[5:0] | rob_valid_35; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10660 = 6'h24 == allocate_ptr[5:0] | rob_valid_36; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10661 = 6'h25 == allocate_ptr[5:0] | rob_valid_37; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10662 = 6'h26 == allocate_ptr[5:0] | rob_valid_38; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10663 = 6'h27 == allocate_ptr[5:0] | rob_valid_39; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10664 = 6'h28 == allocate_ptr[5:0] | rob_valid_40; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10665 = 6'h29 == allocate_ptr[5:0] | rob_valid_41; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10666 = 6'h2a == allocate_ptr[5:0] | rob_valid_42; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10667 = 6'h2b == allocate_ptr[5:0] | rob_valid_43; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10668 = 6'h2c == allocate_ptr[5:0] | rob_valid_44; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10669 = 6'h2d == allocate_ptr[5:0] | rob_valid_45; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10670 = 6'h2e == allocate_ptr[5:0] | rob_valid_46; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10671 = 6'h2f == allocate_ptr[5:0] | rob_valid_47; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10672 = 6'h30 == allocate_ptr[5:0] | rob_valid_48; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10673 = 6'h31 == allocate_ptr[5:0] | rob_valid_49; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10674 = 6'h32 == allocate_ptr[5:0] | rob_valid_50; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10675 = 6'h33 == allocate_ptr[5:0] | rob_valid_51; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10676 = 6'h34 == allocate_ptr[5:0] | rob_valid_52; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10677 = 6'h35 == allocate_ptr[5:0] | rob_valid_53; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10678 = 6'h36 == allocate_ptr[5:0] | rob_valid_54; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10679 = 6'h37 == allocate_ptr[5:0] | rob_valid_55; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10680 = 6'h38 == allocate_ptr[5:0] | rob_valid_56; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10681 = 6'h39 == allocate_ptr[5:0] | rob_valid_57; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10682 = 6'h3a == allocate_ptr[5:0] | rob_valid_58; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10683 = 6'h3b == allocate_ptr[5:0] | rob_valid_59; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10684 = 6'h3c == allocate_ptr[5:0] | rob_valid_60; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10685 = 6'h3d == allocate_ptr[5:0] | rob_valid_61; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10686 = 6'h3e == allocate_ptr[5:0] | rob_valid_62; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10687 = 6'h3f == allocate_ptr[5:0] | rob_valid_63; // @[rob.scala 127:{33,33} 81:28]
  wire  _GEN_10688 = 6'h0 == allocate_ptr[5:0] ? 1'h0 : rob_done_0; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10689 = 6'h1 == allocate_ptr[5:0] ? 1'h0 : rob_done_1; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10690 = 6'h2 == allocate_ptr[5:0] ? 1'h0 : rob_done_2; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10691 = 6'h3 == allocate_ptr[5:0] ? 1'h0 : rob_done_3; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10692 = 6'h4 == allocate_ptr[5:0] ? 1'h0 : rob_done_4; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10693 = 6'h5 == allocate_ptr[5:0] ? 1'h0 : rob_done_5; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10694 = 6'h6 == allocate_ptr[5:0] ? 1'h0 : rob_done_6; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10695 = 6'h7 == allocate_ptr[5:0] ? 1'h0 : rob_done_7; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10696 = 6'h8 == allocate_ptr[5:0] ? 1'h0 : rob_done_8; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10697 = 6'h9 == allocate_ptr[5:0] ? 1'h0 : rob_done_9; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10698 = 6'ha == allocate_ptr[5:0] ? 1'h0 : rob_done_10; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10699 = 6'hb == allocate_ptr[5:0] ? 1'h0 : rob_done_11; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10700 = 6'hc == allocate_ptr[5:0] ? 1'h0 : rob_done_12; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10701 = 6'hd == allocate_ptr[5:0] ? 1'h0 : rob_done_13; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10702 = 6'he == allocate_ptr[5:0] ? 1'h0 : rob_done_14; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10703 = 6'hf == allocate_ptr[5:0] ? 1'h0 : rob_done_15; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10704 = 6'h10 == allocate_ptr[5:0] ? 1'h0 : rob_done_16; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10705 = 6'h11 == allocate_ptr[5:0] ? 1'h0 : rob_done_17; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10706 = 6'h12 == allocate_ptr[5:0] ? 1'h0 : rob_done_18; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10707 = 6'h13 == allocate_ptr[5:0] ? 1'h0 : rob_done_19; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10708 = 6'h14 == allocate_ptr[5:0] ? 1'h0 : rob_done_20; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10709 = 6'h15 == allocate_ptr[5:0] ? 1'h0 : rob_done_21; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10710 = 6'h16 == allocate_ptr[5:0] ? 1'h0 : rob_done_22; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10711 = 6'h17 == allocate_ptr[5:0] ? 1'h0 : rob_done_23; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10712 = 6'h18 == allocate_ptr[5:0] ? 1'h0 : rob_done_24; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10713 = 6'h19 == allocate_ptr[5:0] ? 1'h0 : rob_done_25; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10714 = 6'h1a == allocate_ptr[5:0] ? 1'h0 : rob_done_26; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10715 = 6'h1b == allocate_ptr[5:0] ? 1'h0 : rob_done_27; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10716 = 6'h1c == allocate_ptr[5:0] ? 1'h0 : rob_done_28; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10717 = 6'h1d == allocate_ptr[5:0] ? 1'h0 : rob_done_29; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10718 = 6'h1e == allocate_ptr[5:0] ? 1'h0 : rob_done_30; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10719 = 6'h1f == allocate_ptr[5:0] ? 1'h0 : rob_done_31; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10720 = 6'h20 == allocate_ptr[5:0] ? 1'h0 : rob_done_32; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10721 = 6'h21 == allocate_ptr[5:0] ? 1'h0 : rob_done_33; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10722 = 6'h22 == allocate_ptr[5:0] ? 1'h0 : rob_done_34; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10723 = 6'h23 == allocate_ptr[5:0] ? 1'h0 : rob_done_35; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10724 = 6'h24 == allocate_ptr[5:0] ? 1'h0 : rob_done_36; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10725 = 6'h25 == allocate_ptr[5:0] ? 1'h0 : rob_done_37; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10726 = 6'h26 == allocate_ptr[5:0] ? 1'h0 : rob_done_38; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10727 = 6'h27 == allocate_ptr[5:0] ? 1'h0 : rob_done_39; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10728 = 6'h28 == allocate_ptr[5:0] ? 1'h0 : rob_done_40; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10729 = 6'h29 == allocate_ptr[5:0] ? 1'h0 : rob_done_41; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10730 = 6'h2a == allocate_ptr[5:0] ? 1'h0 : rob_done_42; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10731 = 6'h2b == allocate_ptr[5:0] ? 1'h0 : rob_done_43; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10732 = 6'h2c == allocate_ptr[5:0] ? 1'h0 : rob_done_44; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10733 = 6'h2d == allocate_ptr[5:0] ? 1'h0 : rob_done_45; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10734 = 6'h2e == allocate_ptr[5:0] ? 1'h0 : rob_done_46; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10735 = 6'h2f == allocate_ptr[5:0] ? 1'h0 : rob_done_47; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10736 = 6'h30 == allocate_ptr[5:0] ? 1'h0 : rob_done_48; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10737 = 6'h31 == allocate_ptr[5:0] ? 1'h0 : rob_done_49; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10738 = 6'h32 == allocate_ptr[5:0] ? 1'h0 : rob_done_50; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10739 = 6'h33 == allocate_ptr[5:0] ? 1'h0 : rob_done_51; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10740 = 6'h34 == allocate_ptr[5:0] ? 1'h0 : rob_done_52; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10741 = 6'h35 == allocate_ptr[5:0] ? 1'h0 : rob_done_53; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10742 = 6'h36 == allocate_ptr[5:0] ? 1'h0 : rob_done_54; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10743 = 6'h37 == allocate_ptr[5:0] ? 1'h0 : rob_done_55; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10744 = 6'h38 == allocate_ptr[5:0] ? 1'h0 : rob_done_56; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10745 = 6'h39 == allocate_ptr[5:0] ? 1'h0 : rob_done_57; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10746 = 6'h3a == allocate_ptr[5:0] ? 1'h0 : rob_done_58; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10747 = 6'h3b == allocate_ptr[5:0] ? 1'h0 : rob_done_59; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10748 = 6'h3c == allocate_ptr[5:0] ? 1'h0 : rob_done_60; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10749 = 6'h3d == allocate_ptr[5:0] ? 1'h0 : rob_done_61; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10750 = 6'h3e == allocate_ptr[5:0] ? 1'h0 : rob_done_62; // @[rob.scala 128:{32,32} 84:27]
  wire  _GEN_10751 = 6'h3f == allocate_ptr[5:0] ? 1'h0 : rob_done_63; // @[rob.scala 128:{32,32} 84:27]
  wire [31:0] _GEN_10816 = 6'h0 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8704; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10817 = 6'h1 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8705; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10818 = 6'h2 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8706; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10819 = 6'h3 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8707; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10820 = 6'h4 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8708; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10821 = 6'h5 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8709; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10822 = 6'h6 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8710; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10823 = 6'h7 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8711; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10824 = 6'h8 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8712; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10825 = 6'h9 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8713; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10826 = 6'ha == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8714; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10827 = 6'hb == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8715; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10828 = 6'hc == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8716; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10829 = 6'hd == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8717; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10830 = 6'he == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8718; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10831 = 6'hf == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8719; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10832 = 6'h10 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8720; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10833 = 6'h11 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8721; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10834 = 6'h12 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8722; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10835 = 6'h13 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8723; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10836 = 6'h14 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8724; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10837 = 6'h15 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8725; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10838 = 6'h16 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8726; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10839 = 6'h17 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8727; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10840 = 6'h18 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8728; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10841 = 6'h19 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8729; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10842 = 6'h1a == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8730; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10843 = 6'h1b == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8731; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10844 = 6'h1c == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8732; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10845 = 6'h1d == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8733; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10846 = 6'h1e == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8734; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10847 = 6'h1f == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8735; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10848 = 6'h20 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8736; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10849 = 6'h21 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8737; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10850 = 6'h22 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8738; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10851 = 6'h23 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8739; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10852 = 6'h24 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8740; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10853 = 6'h25 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8741; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10854 = 6'h26 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8742; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10855 = 6'h27 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8743; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10856 = 6'h28 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8744; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10857 = 6'h29 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8745; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10858 = 6'h2a == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8746; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10859 = 6'h2b == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8747; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10860 = 6'h2c == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8748; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10861 = 6'h2d == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8749; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10862 = 6'h2e == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8750; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10863 = 6'h2f == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8751; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10864 = 6'h30 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8752; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10865 = 6'h31 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8753; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10866 = 6'h32 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8754; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10867 = 6'h33 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8755; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10868 = 6'h34 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8756; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10869 = 6'h35 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8757; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10870 = 6'h36 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8758; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10871 = 6'h37 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8759; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10872 = 6'h38 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8760; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10873 = 6'h39 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8761; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10874 = 6'h3a == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8762; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10875 = 6'h3b == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8763; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10876 = 6'h3c == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8764; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10877 = 6'h3d == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8765; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10878 = 6'h3e == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8766; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10879 = 6'h3f == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_pc : _GEN_8767; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10880 = 6'h0 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8768; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10881 = 6'h1 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8769; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10882 = 6'h2 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8770; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10883 = 6'h3 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8771; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10884 = 6'h4 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8772; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10885 = 6'h5 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8773; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10886 = 6'h6 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8774; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10887 = 6'h7 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8775; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10888 = 6'h8 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8776; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10889 = 6'h9 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8777; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10890 = 6'ha == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8778; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10891 = 6'hb == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8779; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10892 = 6'hc == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8780; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10893 = 6'hd == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8781; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10894 = 6'he == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8782; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10895 = 6'hf == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8783; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10896 = 6'h10 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8784; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10897 = 6'h11 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8785; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10898 = 6'h12 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8786; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10899 = 6'h13 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8787; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10900 = 6'h14 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8788; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10901 = 6'h15 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8789; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10902 = 6'h16 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8790; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10903 = 6'h17 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8791; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10904 = 6'h18 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8792; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10905 = 6'h19 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8793; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10906 = 6'h1a == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8794; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10907 = 6'h1b == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8795; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10908 = 6'h1c == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8796; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10909 = 6'h1d == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8797; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10910 = 6'h1e == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8798; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10911 = 6'h1f == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8799; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10912 = 6'h20 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8800; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10913 = 6'h21 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8801; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10914 = 6'h22 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8802; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10915 = 6'h23 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8803; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10916 = 6'h24 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8804; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10917 = 6'h25 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8805; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10918 = 6'h26 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8806; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10919 = 6'h27 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8807; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10920 = 6'h28 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8808; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10921 = 6'h29 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8809; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10922 = 6'h2a == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8810; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10923 = 6'h2b == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8811; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10924 = 6'h2c == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8812; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10925 = 6'h2d == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8813; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10926 = 6'h2e == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8814; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10927 = 6'h2f == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8815; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10928 = 6'h30 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8816; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10929 = 6'h31 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8817; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10930 = 6'h32 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8818; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10931 = 6'h33 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8819; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10932 = 6'h34 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8820; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10933 = 6'h35 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8821; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10934 = 6'h36 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8822; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10935 = 6'h37 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8823; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10936 = 6'h38 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8824; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10937 = 6'h39 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8825; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10938 = 6'h3a == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8826; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10939 = 6'h3b == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8827; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10940 = 6'h3c == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8828; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10941 = 6'h3d == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8829; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10942 = 6'h3e == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8830; // @[rob.scala 129:{35,35}]
  wire [31:0] _GEN_10943 = 6'h3f == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_inst : _GEN_8831; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10944 = 6'h0 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8832; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10945 = 6'h1 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8833; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10946 = 6'h2 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8834; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10947 = 6'h3 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8835; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10948 = 6'h4 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8836; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10949 = 6'h5 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8837; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10950 = 6'h6 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8838; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10951 = 6'h7 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8839; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10952 = 6'h8 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8840; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10953 = 6'h9 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8841; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10954 = 6'ha == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8842; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10955 = 6'hb == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8843; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10956 = 6'hc == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8844; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10957 = 6'hd == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8845; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10958 = 6'he == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8846; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10959 = 6'hf == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8847; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10960 = 6'h10 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8848; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10961 = 6'h11 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8849; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10962 = 6'h12 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8850; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10963 = 6'h13 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8851; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10964 = 6'h14 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8852; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10965 = 6'h15 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8853; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10966 = 6'h16 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8854; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10967 = 6'h17 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8855; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10968 = 6'h18 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8856; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10969 = 6'h19 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8857; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10970 = 6'h1a == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8858; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10971 = 6'h1b == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8859; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10972 = 6'h1c == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8860; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10973 = 6'h1d == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8861; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10974 = 6'h1e == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8862; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10975 = 6'h1f == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8863; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10976 = 6'h20 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8864; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10977 = 6'h21 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8865; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10978 = 6'h22 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8866; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10979 = 6'h23 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8867; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10980 = 6'h24 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8868; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10981 = 6'h25 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8869; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10982 = 6'h26 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8870; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10983 = 6'h27 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8871; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10984 = 6'h28 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8872; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10985 = 6'h29 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8873; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10986 = 6'h2a == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8874; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10987 = 6'h2b == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8875; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10988 = 6'h2c == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8876; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10989 = 6'h2d == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8877; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10990 = 6'h2e == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8878; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10991 = 6'h2f == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8879; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10992 = 6'h30 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8880; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10993 = 6'h31 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8881; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10994 = 6'h32 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8882; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10995 = 6'h33 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8883; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10996 = 6'h34 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8884; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10997 = 6'h35 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8885; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10998 = 6'h36 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8886; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_10999 = 6'h37 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8887; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11000 = 6'h38 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8888; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11001 = 6'h39 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8889; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11002 = 6'h3a == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8890; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11003 = 6'h3b == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8891; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11004 = 6'h3c == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8892; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11005 = 6'h3d == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8893; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11006 = 6'h3e == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8894; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11007 = 6'h3f == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_func_code : _GEN_8895; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11328 = 6'h0 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9216; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11329 = 6'h1 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9217; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11330 = 6'h2 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9218; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11331 = 6'h3 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9219; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11332 = 6'h4 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9220; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11333 = 6'h5 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9221; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11334 = 6'h6 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9222; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11335 = 6'h7 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9223; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11336 = 6'h8 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9224; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11337 = 6'h9 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9225; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11338 = 6'ha == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9226; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11339 = 6'hb == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9227; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11340 = 6'hc == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9228; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11341 = 6'hd == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9229; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11342 = 6'he == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9230; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11343 = 6'hf == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9231; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11344 = 6'h10 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9232; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11345 = 6'h11 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9233; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11346 = 6'h12 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9234; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11347 = 6'h13 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9235; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11348 = 6'h14 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9236; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11349 = 6'h15 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9237; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11350 = 6'h16 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9238; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11351 = 6'h17 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9239; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11352 = 6'h18 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9240; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11353 = 6'h19 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9241; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11354 = 6'h1a == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9242; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11355 = 6'h1b == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9243; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11356 = 6'h1c == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9244; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11357 = 6'h1d == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9245; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11358 = 6'h1e == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9246; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11359 = 6'h1f == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9247; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11360 = 6'h20 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9248; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11361 = 6'h21 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9249; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11362 = 6'h22 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9250; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11363 = 6'h23 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9251; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11364 = 6'h24 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9252; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11365 = 6'h25 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9253; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11366 = 6'h26 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9254; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11367 = 6'h27 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9255; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11368 = 6'h28 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9256; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11369 = 6'h29 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9257; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11370 = 6'h2a == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9258; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11371 = 6'h2b == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9259; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11372 = 6'h2c == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9260; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11373 = 6'h2d == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9261; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11374 = 6'h2e == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9262; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11375 = 6'h2f == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9263; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11376 = 6'h30 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9264; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11377 = 6'h31 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9265; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11378 = 6'h32 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9266; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11379 = 6'h33 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9267; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11380 = 6'h34 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9268; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11381 = 6'h35 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9269; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11382 = 6'h36 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9270; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11383 = 6'h37 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9271; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11384 = 6'h38 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9272; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11385 = 6'h39 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9273; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11386 = 6'h3a == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9274; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11387 = 6'h3b == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9275; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11388 = 6'h3c == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9276; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11389 = 6'h3d == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9277; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11390 = 6'h3e == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9278; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11391 = 6'h3f == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_phy_dst : _GEN_9279; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11392 = 6'h0 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9280; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11393 = 6'h1 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9281; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11394 = 6'h2 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9282; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11395 = 6'h3 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9283; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11396 = 6'h4 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9284; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11397 = 6'h5 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9285; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11398 = 6'h6 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9286; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11399 = 6'h7 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9287; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11400 = 6'h8 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9288; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11401 = 6'h9 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9289; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11402 = 6'ha == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9290; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11403 = 6'hb == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9291; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11404 = 6'hc == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9292; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11405 = 6'hd == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9293; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11406 = 6'he == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9294; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11407 = 6'hf == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9295; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11408 = 6'h10 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9296; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11409 = 6'h11 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9297; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11410 = 6'h12 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9298; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11411 = 6'h13 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9299; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11412 = 6'h14 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9300; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11413 = 6'h15 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9301; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11414 = 6'h16 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9302; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11415 = 6'h17 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9303; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11416 = 6'h18 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9304; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11417 = 6'h19 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9305; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11418 = 6'h1a == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9306; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11419 = 6'h1b == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9307; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11420 = 6'h1c == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9308; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11421 = 6'h1d == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9309; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11422 = 6'h1e == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9310; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11423 = 6'h1f == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9311; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11424 = 6'h20 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9312; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11425 = 6'h21 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9313; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11426 = 6'h22 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9314; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11427 = 6'h23 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9315; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11428 = 6'h24 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9316; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11429 = 6'h25 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9317; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11430 = 6'h26 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9318; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11431 = 6'h27 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9319; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11432 = 6'h28 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9320; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11433 = 6'h29 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9321; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11434 = 6'h2a == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9322; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11435 = 6'h2b == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9323; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11436 = 6'h2c == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9324; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11437 = 6'h2d == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9325; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11438 = 6'h2e == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9326; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11439 = 6'h2f == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9327; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11440 = 6'h30 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9328; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11441 = 6'h31 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9329; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11442 = 6'h32 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9330; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11443 = 6'h33 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9331; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11444 = 6'h34 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9332; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11445 = 6'h35 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9333; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11446 = 6'h36 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9334; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11447 = 6'h37 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9335; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11448 = 6'h38 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9336; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11449 = 6'h39 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9337; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11450 = 6'h3a == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9338; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11451 = 6'h3b == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9339; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11452 = 6'h3c == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9340; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11453 = 6'h3d == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9341; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11454 = 6'h3e == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9342; // @[rob.scala 129:{35,35}]
  wire [6:0] _GEN_11455 = 6'h3f == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_stale_dst : _GEN_9343; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11456 = 6'h0 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9344; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11457 = 6'h1 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9345; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11458 = 6'h2 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9346; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11459 = 6'h3 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9347; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11460 = 6'h4 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9348; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11461 = 6'h5 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9349; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11462 = 6'h6 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9350; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11463 = 6'h7 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9351; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11464 = 6'h8 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9352; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11465 = 6'h9 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9353; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11466 = 6'ha == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9354; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11467 = 6'hb == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9355; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11468 = 6'hc == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9356; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11469 = 6'hd == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9357; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11470 = 6'he == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9358; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11471 = 6'hf == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9359; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11472 = 6'h10 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9360; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11473 = 6'h11 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9361; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11474 = 6'h12 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9362; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11475 = 6'h13 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9363; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11476 = 6'h14 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9364; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11477 = 6'h15 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9365; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11478 = 6'h16 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9366; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11479 = 6'h17 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9367; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11480 = 6'h18 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9368; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11481 = 6'h19 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9369; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11482 = 6'h1a == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9370; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11483 = 6'h1b == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9371; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11484 = 6'h1c == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9372; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11485 = 6'h1d == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9373; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11486 = 6'h1e == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9374; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11487 = 6'h1f == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9375; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11488 = 6'h20 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9376; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11489 = 6'h21 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9377; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11490 = 6'h22 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9378; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11491 = 6'h23 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9379; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11492 = 6'h24 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9380; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11493 = 6'h25 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9381; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11494 = 6'h26 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9382; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11495 = 6'h27 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9383; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11496 = 6'h28 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9384; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11497 = 6'h29 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9385; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11498 = 6'h2a == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9386; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11499 = 6'h2b == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9387; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11500 = 6'h2c == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9388; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11501 = 6'h2d == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9389; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11502 = 6'h2e == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9390; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11503 = 6'h2f == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9391; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11504 = 6'h30 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9392; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11505 = 6'h31 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9393; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11506 = 6'h32 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9394; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11507 = 6'h33 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9395; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11508 = 6'h34 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9396; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11509 = 6'h35 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9397; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11510 = 6'h36 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9398; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11511 = 6'h37 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9399; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11512 = 6'h38 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9400; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11513 = 6'h39 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9401; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11514 = 6'h3a == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9402; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11515 = 6'h3b == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9403; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11516 = 6'h3c == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9404; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11517 = 6'h3d == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9405; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11518 = 6'h3e == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9406; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_11519 = 6'h3f == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_arch_dst : _GEN_9407; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12160 = 6'h0 == _is_full_T_4[5:0] ? 64'h0 : _GEN_10048; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12161 = 6'h1 == _is_full_T_4[5:0] ? 64'h0 : _GEN_10049; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12162 = 6'h2 == _is_full_T_4[5:0] ? 64'h0 : _GEN_10050; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12163 = 6'h3 == _is_full_T_4[5:0] ? 64'h0 : _GEN_10051; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12164 = 6'h4 == _is_full_T_4[5:0] ? 64'h0 : _GEN_10052; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12165 = 6'h5 == _is_full_T_4[5:0] ? 64'h0 : _GEN_10053; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12166 = 6'h6 == _is_full_T_4[5:0] ? 64'h0 : _GEN_10054; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12167 = 6'h7 == _is_full_T_4[5:0] ? 64'h0 : _GEN_10055; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12168 = 6'h8 == _is_full_T_4[5:0] ? 64'h0 : _GEN_10056; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12169 = 6'h9 == _is_full_T_4[5:0] ? 64'h0 : _GEN_10057; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12170 = 6'ha == _is_full_T_4[5:0] ? 64'h0 : _GEN_10058; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12171 = 6'hb == _is_full_T_4[5:0] ? 64'h0 : _GEN_10059; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12172 = 6'hc == _is_full_T_4[5:0] ? 64'h0 : _GEN_10060; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12173 = 6'hd == _is_full_T_4[5:0] ? 64'h0 : _GEN_10061; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12174 = 6'he == _is_full_T_4[5:0] ? 64'h0 : _GEN_10062; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12175 = 6'hf == _is_full_T_4[5:0] ? 64'h0 : _GEN_10063; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12176 = 6'h10 == _is_full_T_4[5:0] ? 64'h0 : _GEN_10064; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12177 = 6'h11 == _is_full_T_4[5:0] ? 64'h0 : _GEN_10065; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12178 = 6'h12 == _is_full_T_4[5:0] ? 64'h0 : _GEN_10066; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12179 = 6'h13 == _is_full_T_4[5:0] ? 64'h0 : _GEN_10067; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12180 = 6'h14 == _is_full_T_4[5:0] ? 64'h0 : _GEN_10068; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12181 = 6'h15 == _is_full_T_4[5:0] ? 64'h0 : _GEN_10069; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12182 = 6'h16 == _is_full_T_4[5:0] ? 64'h0 : _GEN_10070; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12183 = 6'h17 == _is_full_T_4[5:0] ? 64'h0 : _GEN_10071; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12184 = 6'h18 == _is_full_T_4[5:0] ? 64'h0 : _GEN_10072; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12185 = 6'h19 == _is_full_T_4[5:0] ? 64'h0 : _GEN_10073; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12186 = 6'h1a == _is_full_T_4[5:0] ? 64'h0 : _GEN_10074; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12187 = 6'h1b == _is_full_T_4[5:0] ? 64'h0 : _GEN_10075; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12188 = 6'h1c == _is_full_T_4[5:0] ? 64'h0 : _GEN_10076; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12189 = 6'h1d == _is_full_T_4[5:0] ? 64'h0 : _GEN_10077; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12190 = 6'h1e == _is_full_T_4[5:0] ? 64'h0 : _GEN_10078; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12191 = 6'h1f == _is_full_T_4[5:0] ? 64'h0 : _GEN_10079; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12192 = 6'h20 == _is_full_T_4[5:0] ? 64'h0 : _GEN_10080; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12193 = 6'h21 == _is_full_T_4[5:0] ? 64'h0 : _GEN_10081; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12194 = 6'h22 == _is_full_T_4[5:0] ? 64'h0 : _GEN_10082; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12195 = 6'h23 == _is_full_T_4[5:0] ? 64'h0 : _GEN_10083; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12196 = 6'h24 == _is_full_T_4[5:0] ? 64'h0 : _GEN_10084; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12197 = 6'h25 == _is_full_T_4[5:0] ? 64'h0 : _GEN_10085; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12198 = 6'h26 == _is_full_T_4[5:0] ? 64'h0 : _GEN_10086; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12199 = 6'h27 == _is_full_T_4[5:0] ? 64'h0 : _GEN_10087; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12200 = 6'h28 == _is_full_T_4[5:0] ? 64'h0 : _GEN_10088; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12201 = 6'h29 == _is_full_T_4[5:0] ? 64'h0 : _GEN_10089; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12202 = 6'h2a == _is_full_T_4[5:0] ? 64'h0 : _GEN_10090; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12203 = 6'h2b == _is_full_T_4[5:0] ? 64'h0 : _GEN_10091; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12204 = 6'h2c == _is_full_T_4[5:0] ? 64'h0 : _GEN_10092; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12205 = 6'h2d == _is_full_T_4[5:0] ? 64'h0 : _GEN_10093; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12206 = 6'h2e == _is_full_T_4[5:0] ? 64'h0 : _GEN_10094; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12207 = 6'h2f == _is_full_T_4[5:0] ? 64'h0 : _GEN_10095; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12208 = 6'h30 == _is_full_T_4[5:0] ? 64'h0 : _GEN_10096; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12209 = 6'h31 == _is_full_T_4[5:0] ? 64'h0 : _GEN_10097; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12210 = 6'h32 == _is_full_T_4[5:0] ? 64'h0 : _GEN_10098; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12211 = 6'h33 == _is_full_T_4[5:0] ? 64'h0 : _GEN_10099; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12212 = 6'h34 == _is_full_T_4[5:0] ? 64'h0 : _GEN_10100; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12213 = 6'h35 == _is_full_T_4[5:0] ? 64'h0 : _GEN_10101; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12214 = 6'h36 == _is_full_T_4[5:0] ? 64'h0 : _GEN_10102; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12215 = 6'h37 == _is_full_T_4[5:0] ? 64'h0 : _GEN_10103; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12216 = 6'h38 == _is_full_T_4[5:0] ? 64'h0 : _GEN_10104; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12217 = 6'h39 == _is_full_T_4[5:0] ? 64'h0 : _GEN_10105; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12218 = 6'h3a == _is_full_T_4[5:0] ? 64'h0 : _GEN_10106; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12219 = 6'h3b == _is_full_T_4[5:0] ? 64'h0 : _GEN_10107; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12220 = 6'h3c == _is_full_T_4[5:0] ? 64'h0 : _GEN_10108; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12221 = 6'h3d == _is_full_T_4[5:0] ? 64'h0 : _GEN_10109; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12222 = 6'h3e == _is_full_T_4[5:0] ? 64'h0 : _GEN_10110; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12223 = 6'h3f == _is_full_T_4[5:0] ? 64'h0 : _GEN_10111; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12224 = 6'h0 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10112; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12225 = 6'h1 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10113; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12226 = 6'h2 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10114; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12227 = 6'h3 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10115; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12228 = 6'h4 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10116; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12229 = 6'h5 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10117; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12230 = 6'h6 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10118; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12231 = 6'h7 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10119; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12232 = 6'h8 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10120; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12233 = 6'h9 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10121; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12234 = 6'ha == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10122; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12235 = 6'hb == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10123; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12236 = 6'hc == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10124; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12237 = 6'hd == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10125; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12238 = 6'he == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10126; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12239 = 6'hf == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10127; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12240 = 6'h10 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10128; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12241 = 6'h11 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10129; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12242 = 6'h12 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10130; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12243 = 6'h13 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10131; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12244 = 6'h14 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10132; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12245 = 6'h15 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10133; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12246 = 6'h16 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10134; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12247 = 6'h17 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10135; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12248 = 6'h18 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10136; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12249 = 6'h19 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10137; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12250 = 6'h1a == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10138; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12251 = 6'h1b == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10139; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12252 = 6'h1c == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10140; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12253 = 6'h1d == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10141; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12254 = 6'h1e == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10142; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12255 = 6'h1f == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10143; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12256 = 6'h20 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10144; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12257 = 6'h21 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10145; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12258 = 6'h22 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10146; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12259 = 6'h23 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10147; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12260 = 6'h24 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10148; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12261 = 6'h25 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10149; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12262 = 6'h26 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10150; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12263 = 6'h27 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10151; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12264 = 6'h28 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10152; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12265 = 6'h29 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10153; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12266 = 6'h2a == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10154; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12267 = 6'h2b == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10155; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12268 = 6'h2c == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10156; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12269 = 6'h2d == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10157; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12270 = 6'h2e == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10158; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12271 = 6'h2f == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10159; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12272 = 6'h30 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10160; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12273 = 6'h31 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10161; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12274 = 6'h32 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10162; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12275 = 6'h33 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10163; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12276 = 6'h34 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10164; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12277 = 6'h35 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10165; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12278 = 6'h36 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10166; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12279 = 6'h37 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10167; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12280 = 6'h38 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10168; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12281 = 6'h39 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10169; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12282 = 6'h3a == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10170; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12283 = 6'h3b == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10171; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12284 = 6'h3c == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10172; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12285 = 6'h3d == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10173; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12286 = 6'h3e == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10174; // @[rob.scala 129:{35,35}]
  wire [63:0] _GEN_12287 = 6'h3f == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_src1_value : _GEN_10175; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12544 = 6'h0 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10432; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12545 = 6'h1 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10433; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12546 = 6'h2 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10434; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12547 = 6'h3 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10435; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12548 = 6'h4 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10436; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12549 = 6'h5 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10437; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12550 = 6'h6 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10438; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12551 = 6'h7 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10439; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12552 = 6'h8 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10440; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12553 = 6'h9 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10441; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12554 = 6'ha == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10442; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12555 = 6'hb == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10443; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12556 = 6'hc == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10444; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12557 = 6'hd == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10445; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12558 = 6'he == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10446; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12559 = 6'hf == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10447; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12560 = 6'h10 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10448; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12561 = 6'h11 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10449; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12562 = 6'h12 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10450; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12563 = 6'h13 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10451; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12564 = 6'h14 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10452; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12565 = 6'h15 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10453; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12566 = 6'h16 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10454; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12567 = 6'h17 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10455; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12568 = 6'h18 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10456; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12569 = 6'h19 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10457; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12570 = 6'h1a == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10458; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12571 = 6'h1b == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10459; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12572 = 6'h1c == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10460; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12573 = 6'h1d == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10461; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12574 = 6'h1e == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10462; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12575 = 6'h1f == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10463; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12576 = 6'h20 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10464; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12577 = 6'h21 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10465; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12578 = 6'h22 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10466; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12579 = 6'h23 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10467; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12580 = 6'h24 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10468; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12581 = 6'h25 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10469; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12582 = 6'h26 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10470; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12583 = 6'h27 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10471; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12584 = 6'h28 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10472; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12585 = 6'h29 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10473; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12586 = 6'h2a == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10474; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12587 = 6'h2b == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10475; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12588 = 6'h2c == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10476; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12589 = 6'h2d == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10477; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12590 = 6'h2e == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10478; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12591 = 6'h2f == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10479; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12592 = 6'h30 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10480; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12593 = 6'h31 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10481; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12594 = 6'h32 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10482; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12595 = 6'h33 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10483; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12596 = 6'h34 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10484; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12597 = 6'h35 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10485; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12598 = 6'h36 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10486; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12599 = 6'h37 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10487; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12600 = 6'h38 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10488; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12601 = 6'h39 == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10489; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12602 = 6'h3a == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10490; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12603 = 6'h3b == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10491; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12604 = 6'h3c == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10492; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12605 = 6'h3d == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10493; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12606 = 6'h3e == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10494; // @[rob.scala 129:{35,35}]
  wire [4:0] _GEN_12607 = 6'h3f == _is_full_T_4[5:0] ? io_i_rob_allocation_reqs_1_uop_alu_sel : _GEN_10495; // @[rob.scala 129:{35,35}]
  wire  _GEN_12736 = 6'h0 == _is_full_T_4[5:0] | _GEN_10624; // @[rob.scala 130:{37,37}]
  wire  _GEN_12737 = 6'h1 == _is_full_T_4[5:0] | _GEN_10625; // @[rob.scala 130:{37,37}]
  wire  _GEN_12738 = 6'h2 == _is_full_T_4[5:0] | _GEN_10626; // @[rob.scala 130:{37,37}]
  wire  _GEN_12739 = 6'h3 == _is_full_T_4[5:0] | _GEN_10627; // @[rob.scala 130:{37,37}]
  wire  _GEN_12740 = 6'h4 == _is_full_T_4[5:0] | _GEN_10628; // @[rob.scala 130:{37,37}]
  wire  _GEN_12741 = 6'h5 == _is_full_T_4[5:0] | _GEN_10629; // @[rob.scala 130:{37,37}]
  wire  _GEN_12742 = 6'h6 == _is_full_T_4[5:0] | _GEN_10630; // @[rob.scala 130:{37,37}]
  wire  _GEN_12743 = 6'h7 == _is_full_T_4[5:0] | _GEN_10631; // @[rob.scala 130:{37,37}]
  wire  _GEN_12744 = 6'h8 == _is_full_T_4[5:0] | _GEN_10632; // @[rob.scala 130:{37,37}]
  wire  _GEN_12745 = 6'h9 == _is_full_T_4[5:0] | _GEN_10633; // @[rob.scala 130:{37,37}]
  wire  _GEN_12746 = 6'ha == _is_full_T_4[5:0] | _GEN_10634; // @[rob.scala 130:{37,37}]
  wire  _GEN_12747 = 6'hb == _is_full_T_4[5:0] | _GEN_10635; // @[rob.scala 130:{37,37}]
  wire  _GEN_12748 = 6'hc == _is_full_T_4[5:0] | _GEN_10636; // @[rob.scala 130:{37,37}]
  wire  _GEN_12749 = 6'hd == _is_full_T_4[5:0] | _GEN_10637; // @[rob.scala 130:{37,37}]
  wire  _GEN_12750 = 6'he == _is_full_T_4[5:0] | _GEN_10638; // @[rob.scala 130:{37,37}]
  wire  _GEN_12751 = 6'hf == _is_full_T_4[5:0] | _GEN_10639; // @[rob.scala 130:{37,37}]
  wire  _GEN_12752 = 6'h10 == _is_full_T_4[5:0] | _GEN_10640; // @[rob.scala 130:{37,37}]
  wire  _GEN_12753 = 6'h11 == _is_full_T_4[5:0] | _GEN_10641; // @[rob.scala 130:{37,37}]
  wire  _GEN_12754 = 6'h12 == _is_full_T_4[5:0] | _GEN_10642; // @[rob.scala 130:{37,37}]
  wire  _GEN_12755 = 6'h13 == _is_full_T_4[5:0] | _GEN_10643; // @[rob.scala 130:{37,37}]
  wire  _GEN_12756 = 6'h14 == _is_full_T_4[5:0] | _GEN_10644; // @[rob.scala 130:{37,37}]
  wire  _GEN_12757 = 6'h15 == _is_full_T_4[5:0] | _GEN_10645; // @[rob.scala 130:{37,37}]
  wire  _GEN_12758 = 6'h16 == _is_full_T_4[5:0] | _GEN_10646; // @[rob.scala 130:{37,37}]
  wire  _GEN_12759 = 6'h17 == _is_full_T_4[5:0] | _GEN_10647; // @[rob.scala 130:{37,37}]
  wire  _GEN_12760 = 6'h18 == _is_full_T_4[5:0] | _GEN_10648; // @[rob.scala 130:{37,37}]
  wire  _GEN_12761 = 6'h19 == _is_full_T_4[5:0] | _GEN_10649; // @[rob.scala 130:{37,37}]
  wire  _GEN_12762 = 6'h1a == _is_full_T_4[5:0] | _GEN_10650; // @[rob.scala 130:{37,37}]
  wire  _GEN_12763 = 6'h1b == _is_full_T_4[5:0] | _GEN_10651; // @[rob.scala 130:{37,37}]
  wire  _GEN_12764 = 6'h1c == _is_full_T_4[5:0] | _GEN_10652; // @[rob.scala 130:{37,37}]
  wire  _GEN_12765 = 6'h1d == _is_full_T_4[5:0] | _GEN_10653; // @[rob.scala 130:{37,37}]
  wire  _GEN_12766 = 6'h1e == _is_full_T_4[5:0] | _GEN_10654; // @[rob.scala 130:{37,37}]
  wire  _GEN_12767 = 6'h1f == _is_full_T_4[5:0] | _GEN_10655; // @[rob.scala 130:{37,37}]
  wire  _GEN_12768 = 6'h20 == _is_full_T_4[5:0] | _GEN_10656; // @[rob.scala 130:{37,37}]
  wire  _GEN_12769 = 6'h21 == _is_full_T_4[5:0] | _GEN_10657; // @[rob.scala 130:{37,37}]
  wire  _GEN_12770 = 6'h22 == _is_full_T_4[5:0] | _GEN_10658; // @[rob.scala 130:{37,37}]
  wire  _GEN_12771 = 6'h23 == _is_full_T_4[5:0] | _GEN_10659; // @[rob.scala 130:{37,37}]
  wire  _GEN_12772 = 6'h24 == _is_full_T_4[5:0] | _GEN_10660; // @[rob.scala 130:{37,37}]
  wire  _GEN_12773 = 6'h25 == _is_full_T_4[5:0] | _GEN_10661; // @[rob.scala 130:{37,37}]
  wire  _GEN_12774 = 6'h26 == _is_full_T_4[5:0] | _GEN_10662; // @[rob.scala 130:{37,37}]
  wire  _GEN_12775 = 6'h27 == _is_full_T_4[5:0] | _GEN_10663; // @[rob.scala 130:{37,37}]
  wire  _GEN_12776 = 6'h28 == _is_full_T_4[5:0] | _GEN_10664; // @[rob.scala 130:{37,37}]
  wire  _GEN_12777 = 6'h29 == _is_full_T_4[5:0] | _GEN_10665; // @[rob.scala 130:{37,37}]
  wire  _GEN_12778 = 6'h2a == _is_full_T_4[5:0] | _GEN_10666; // @[rob.scala 130:{37,37}]
  wire  _GEN_12779 = 6'h2b == _is_full_T_4[5:0] | _GEN_10667; // @[rob.scala 130:{37,37}]
  wire  _GEN_12780 = 6'h2c == _is_full_T_4[5:0] | _GEN_10668; // @[rob.scala 130:{37,37}]
  wire  _GEN_12781 = 6'h2d == _is_full_T_4[5:0] | _GEN_10669; // @[rob.scala 130:{37,37}]
  wire  _GEN_12782 = 6'h2e == _is_full_T_4[5:0] | _GEN_10670; // @[rob.scala 130:{37,37}]
  wire  _GEN_12783 = 6'h2f == _is_full_T_4[5:0] | _GEN_10671; // @[rob.scala 130:{37,37}]
  wire  _GEN_12784 = 6'h30 == _is_full_T_4[5:0] | _GEN_10672; // @[rob.scala 130:{37,37}]
  wire  _GEN_12785 = 6'h31 == _is_full_T_4[5:0] | _GEN_10673; // @[rob.scala 130:{37,37}]
  wire  _GEN_12786 = 6'h32 == _is_full_T_4[5:0] | _GEN_10674; // @[rob.scala 130:{37,37}]
  wire  _GEN_12787 = 6'h33 == _is_full_T_4[5:0] | _GEN_10675; // @[rob.scala 130:{37,37}]
  wire  _GEN_12788 = 6'h34 == _is_full_T_4[5:0] | _GEN_10676; // @[rob.scala 130:{37,37}]
  wire  _GEN_12789 = 6'h35 == _is_full_T_4[5:0] | _GEN_10677; // @[rob.scala 130:{37,37}]
  wire  _GEN_12790 = 6'h36 == _is_full_T_4[5:0] | _GEN_10678; // @[rob.scala 130:{37,37}]
  wire  _GEN_12791 = 6'h37 == _is_full_T_4[5:0] | _GEN_10679; // @[rob.scala 130:{37,37}]
  wire  _GEN_12792 = 6'h38 == _is_full_T_4[5:0] | _GEN_10680; // @[rob.scala 130:{37,37}]
  wire  _GEN_12793 = 6'h39 == _is_full_T_4[5:0] | _GEN_10681; // @[rob.scala 130:{37,37}]
  wire  _GEN_12794 = 6'h3a == _is_full_T_4[5:0] | _GEN_10682; // @[rob.scala 130:{37,37}]
  wire  _GEN_12795 = 6'h3b == _is_full_T_4[5:0] | _GEN_10683; // @[rob.scala 130:{37,37}]
  wire  _GEN_12796 = 6'h3c == _is_full_T_4[5:0] | _GEN_10684; // @[rob.scala 130:{37,37}]
  wire  _GEN_12797 = 6'h3d == _is_full_T_4[5:0] | _GEN_10685; // @[rob.scala 130:{37,37}]
  wire  _GEN_12798 = 6'h3e == _is_full_T_4[5:0] | _GEN_10686; // @[rob.scala 130:{37,37}]
  wire  _GEN_12799 = 6'h3f == _is_full_T_4[5:0] | _GEN_10687; // @[rob.scala 130:{37,37}]
  wire  _GEN_12800 = 6'h0 == _is_full_T_4[5:0] ? 1'h0 : _GEN_10688; // @[rob.scala 131:{36,36}]
  wire  _GEN_12801 = 6'h1 == _is_full_T_4[5:0] ? 1'h0 : _GEN_10689; // @[rob.scala 131:{36,36}]
  wire  _GEN_12802 = 6'h2 == _is_full_T_4[5:0] ? 1'h0 : _GEN_10690; // @[rob.scala 131:{36,36}]
  wire  _GEN_12803 = 6'h3 == _is_full_T_4[5:0] ? 1'h0 : _GEN_10691; // @[rob.scala 131:{36,36}]
  wire  _GEN_12804 = 6'h4 == _is_full_T_4[5:0] ? 1'h0 : _GEN_10692; // @[rob.scala 131:{36,36}]
  wire  _GEN_12805 = 6'h5 == _is_full_T_4[5:0] ? 1'h0 : _GEN_10693; // @[rob.scala 131:{36,36}]
  wire  _GEN_12806 = 6'h6 == _is_full_T_4[5:0] ? 1'h0 : _GEN_10694; // @[rob.scala 131:{36,36}]
  wire  _GEN_12807 = 6'h7 == _is_full_T_4[5:0] ? 1'h0 : _GEN_10695; // @[rob.scala 131:{36,36}]
  wire  _GEN_12808 = 6'h8 == _is_full_T_4[5:0] ? 1'h0 : _GEN_10696; // @[rob.scala 131:{36,36}]
  wire  _GEN_12809 = 6'h9 == _is_full_T_4[5:0] ? 1'h0 : _GEN_10697; // @[rob.scala 131:{36,36}]
  wire  _GEN_12810 = 6'ha == _is_full_T_4[5:0] ? 1'h0 : _GEN_10698; // @[rob.scala 131:{36,36}]
  wire  _GEN_12811 = 6'hb == _is_full_T_4[5:0] ? 1'h0 : _GEN_10699; // @[rob.scala 131:{36,36}]
  wire  _GEN_12812 = 6'hc == _is_full_T_4[5:0] ? 1'h0 : _GEN_10700; // @[rob.scala 131:{36,36}]
  wire  _GEN_12813 = 6'hd == _is_full_T_4[5:0] ? 1'h0 : _GEN_10701; // @[rob.scala 131:{36,36}]
  wire  _GEN_12814 = 6'he == _is_full_T_4[5:0] ? 1'h0 : _GEN_10702; // @[rob.scala 131:{36,36}]
  wire  _GEN_12815 = 6'hf == _is_full_T_4[5:0] ? 1'h0 : _GEN_10703; // @[rob.scala 131:{36,36}]
  wire  _GEN_12816 = 6'h10 == _is_full_T_4[5:0] ? 1'h0 : _GEN_10704; // @[rob.scala 131:{36,36}]
  wire  _GEN_12817 = 6'h11 == _is_full_T_4[5:0] ? 1'h0 : _GEN_10705; // @[rob.scala 131:{36,36}]
  wire  _GEN_12818 = 6'h12 == _is_full_T_4[5:0] ? 1'h0 : _GEN_10706; // @[rob.scala 131:{36,36}]
  wire  _GEN_12819 = 6'h13 == _is_full_T_4[5:0] ? 1'h0 : _GEN_10707; // @[rob.scala 131:{36,36}]
  wire  _GEN_12820 = 6'h14 == _is_full_T_4[5:0] ? 1'h0 : _GEN_10708; // @[rob.scala 131:{36,36}]
  wire  _GEN_12821 = 6'h15 == _is_full_T_4[5:0] ? 1'h0 : _GEN_10709; // @[rob.scala 131:{36,36}]
  wire  _GEN_12822 = 6'h16 == _is_full_T_4[5:0] ? 1'h0 : _GEN_10710; // @[rob.scala 131:{36,36}]
  wire  _GEN_12823 = 6'h17 == _is_full_T_4[5:0] ? 1'h0 : _GEN_10711; // @[rob.scala 131:{36,36}]
  wire  _GEN_12824 = 6'h18 == _is_full_T_4[5:0] ? 1'h0 : _GEN_10712; // @[rob.scala 131:{36,36}]
  wire  _GEN_12825 = 6'h19 == _is_full_T_4[5:0] ? 1'h0 : _GEN_10713; // @[rob.scala 131:{36,36}]
  wire  _GEN_12826 = 6'h1a == _is_full_T_4[5:0] ? 1'h0 : _GEN_10714; // @[rob.scala 131:{36,36}]
  wire  _GEN_12827 = 6'h1b == _is_full_T_4[5:0] ? 1'h0 : _GEN_10715; // @[rob.scala 131:{36,36}]
  wire  _GEN_12828 = 6'h1c == _is_full_T_4[5:0] ? 1'h0 : _GEN_10716; // @[rob.scala 131:{36,36}]
  wire  _GEN_12829 = 6'h1d == _is_full_T_4[5:0] ? 1'h0 : _GEN_10717; // @[rob.scala 131:{36,36}]
  wire  _GEN_12830 = 6'h1e == _is_full_T_4[5:0] ? 1'h0 : _GEN_10718; // @[rob.scala 131:{36,36}]
  wire  _GEN_12831 = 6'h1f == _is_full_T_4[5:0] ? 1'h0 : _GEN_10719; // @[rob.scala 131:{36,36}]
  wire  _GEN_12832 = 6'h20 == _is_full_T_4[5:0] ? 1'h0 : _GEN_10720; // @[rob.scala 131:{36,36}]
  wire  _GEN_12833 = 6'h21 == _is_full_T_4[5:0] ? 1'h0 : _GEN_10721; // @[rob.scala 131:{36,36}]
  wire  _GEN_12834 = 6'h22 == _is_full_T_4[5:0] ? 1'h0 : _GEN_10722; // @[rob.scala 131:{36,36}]
  wire  _GEN_12835 = 6'h23 == _is_full_T_4[5:0] ? 1'h0 : _GEN_10723; // @[rob.scala 131:{36,36}]
  wire  _GEN_12836 = 6'h24 == _is_full_T_4[5:0] ? 1'h0 : _GEN_10724; // @[rob.scala 131:{36,36}]
  wire  _GEN_12837 = 6'h25 == _is_full_T_4[5:0] ? 1'h0 : _GEN_10725; // @[rob.scala 131:{36,36}]
  wire  _GEN_12838 = 6'h26 == _is_full_T_4[5:0] ? 1'h0 : _GEN_10726; // @[rob.scala 131:{36,36}]
  wire  _GEN_12839 = 6'h27 == _is_full_T_4[5:0] ? 1'h0 : _GEN_10727; // @[rob.scala 131:{36,36}]
  wire  _GEN_12840 = 6'h28 == _is_full_T_4[5:0] ? 1'h0 : _GEN_10728; // @[rob.scala 131:{36,36}]
  wire  _GEN_12841 = 6'h29 == _is_full_T_4[5:0] ? 1'h0 : _GEN_10729; // @[rob.scala 131:{36,36}]
  wire  _GEN_12842 = 6'h2a == _is_full_T_4[5:0] ? 1'h0 : _GEN_10730; // @[rob.scala 131:{36,36}]
  wire  _GEN_12843 = 6'h2b == _is_full_T_4[5:0] ? 1'h0 : _GEN_10731; // @[rob.scala 131:{36,36}]
  wire  _GEN_12844 = 6'h2c == _is_full_T_4[5:0] ? 1'h0 : _GEN_10732; // @[rob.scala 131:{36,36}]
  wire  _GEN_12845 = 6'h2d == _is_full_T_4[5:0] ? 1'h0 : _GEN_10733; // @[rob.scala 131:{36,36}]
  wire  _GEN_12846 = 6'h2e == _is_full_T_4[5:0] ? 1'h0 : _GEN_10734; // @[rob.scala 131:{36,36}]
  wire  _GEN_12847 = 6'h2f == _is_full_T_4[5:0] ? 1'h0 : _GEN_10735; // @[rob.scala 131:{36,36}]
  wire  _GEN_12848 = 6'h30 == _is_full_T_4[5:0] ? 1'h0 : _GEN_10736; // @[rob.scala 131:{36,36}]
  wire  _GEN_12849 = 6'h31 == _is_full_T_4[5:0] ? 1'h0 : _GEN_10737; // @[rob.scala 131:{36,36}]
  wire  _GEN_12850 = 6'h32 == _is_full_T_4[5:0] ? 1'h0 : _GEN_10738; // @[rob.scala 131:{36,36}]
  wire  _GEN_12851 = 6'h33 == _is_full_T_4[5:0] ? 1'h0 : _GEN_10739; // @[rob.scala 131:{36,36}]
  wire  _GEN_12852 = 6'h34 == _is_full_T_4[5:0] ? 1'h0 : _GEN_10740; // @[rob.scala 131:{36,36}]
  wire  _GEN_12853 = 6'h35 == _is_full_T_4[5:0] ? 1'h0 : _GEN_10741; // @[rob.scala 131:{36,36}]
  wire  _GEN_12854 = 6'h36 == _is_full_T_4[5:0] ? 1'h0 : _GEN_10742; // @[rob.scala 131:{36,36}]
  wire  _GEN_12855 = 6'h37 == _is_full_T_4[5:0] ? 1'h0 : _GEN_10743; // @[rob.scala 131:{36,36}]
  wire  _GEN_12856 = 6'h38 == _is_full_T_4[5:0] ? 1'h0 : _GEN_10744; // @[rob.scala 131:{36,36}]
  wire  _GEN_12857 = 6'h39 == _is_full_T_4[5:0] ? 1'h0 : _GEN_10745; // @[rob.scala 131:{36,36}]
  wire  _GEN_12858 = 6'h3a == _is_full_T_4[5:0] ? 1'h0 : _GEN_10746; // @[rob.scala 131:{36,36}]
  wire  _GEN_12859 = 6'h3b == _is_full_T_4[5:0] ? 1'h0 : _GEN_10747; // @[rob.scala 131:{36,36}]
  wire  _GEN_12860 = 6'h3c == _is_full_T_4[5:0] ? 1'h0 : _GEN_10748; // @[rob.scala 131:{36,36}]
  wire  _GEN_12861 = 6'h3d == _is_full_T_4[5:0] ? 1'h0 : _GEN_10749; // @[rob.scala 131:{36,36}]
  wire  _GEN_12862 = 6'h3e == _is_full_T_4[5:0] ? 1'h0 : _GEN_10750; // @[rob.scala 131:{36,36}]
  wire  _GEN_12863 = 6'h3f == _is_full_T_4[5:0] ? 1'h0 : _GEN_10751; // @[rob.scala 131:{36,36}]
  wire [31:0] _rob_uop_T_pc = io_i_rob_allocation_reqs_0_valid ? io_i_rob_allocation_reqs_0_uop_pc :
    io_i_rob_allocation_reqs_1_uop_pc; // @[rob.scala 134:37]
  wire [31:0] _rob_uop_T_inst = io_i_rob_allocation_reqs_0_valid ? io_i_rob_allocation_reqs_0_uop_inst :
    io_i_rob_allocation_reqs_1_uop_inst; // @[rob.scala 134:37]
  wire [6:0] _rob_uop_T_func_code = io_i_rob_allocation_reqs_0_valid ? io_i_rob_allocation_reqs_0_uop_func_code :
    io_i_rob_allocation_reqs_1_uop_func_code; // @[rob.scala 134:37]
  wire [6:0] _rob_uop_T_phy_dst = io_i_rob_allocation_reqs_0_valid ? io_i_rob_allocation_reqs_0_uop_phy_dst :
    io_i_rob_allocation_reqs_1_uop_phy_dst; // @[rob.scala 134:37]
  wire [6:0] _rob_uop_T_stale_dst = io_i_rob_allocation_reqs_0_valid ? io_i_rob_allocation_reqs_0_uop_stale_dst :
    io_i_rob_allocation_reqs_1_uop_stale_dst; // @[rob.scala 134:37]
  wire [4:0] _rob_uop_T_arch_dst = io_i_rob_allocation_reqs_0_valid ? io_i_rob_allocation_reqs_0_uop_arch_dst :
    io_i_rob_allocation_reqs_1_uop_arch_dst; // @[rob.scala 134:37]
  wire [63:0] _rob_uop_T_src1_value = io_i_rob_allocation_reqs_0_valid ? io_i_rob_allocation_reqs_0_uop_src1_value :
    io_i_rob_allocation_reqs_1_uop_src1_value; // @[rob.scala 134:37]
  wire [4:0] _rob_uop_T_alu_sel = io_i_rob_allocation_reqs_0_valid ? io_i_rob_allocation_reqs_0_uop_alu_sel :
    io_i_rob_allocation_reqs_1_uop_alu_sel; // @[rob.scala 134:37]
  wire [31:0] _GEN_12928 = 6'h0 == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_0_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12929 = 6'h1 == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_1_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12930 = 6'h2 == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_2_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12931 = 6'h3 == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_3_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12932 = 6'h4 == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_4_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12933 = 6'h5 == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_5_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12934 = 6'h6 == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_6_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12935 = 6'h7 == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_7_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12936 = 6'h8 == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_8_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12937 = 6'h9 == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_9_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12938 = 6'ha == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_10_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12939 = 6'hb == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_11_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12940 = 6'hc == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_12_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12941 = 6'hd == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_13_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12942 = 6'he == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_14_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12943 = 6'hf == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_15_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12944 = 6'h10 == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_16_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12945 = 6'h11 == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_17_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12946 = 6'h12 == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_18_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12947 = 6'h13 == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_19_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12948 = 6'h14 == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_20_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12949 = 6'h15 == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_21_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12950 = 6'h16 == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_22_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12951 = 6'h17 == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_23_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12952 = 6'h18 == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_24_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12953 = 6'h19 == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_25_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12954 = 6'h1a == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_26_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12955 = 6'h1b == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_27_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12956 = 6'h1c == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_28_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12957 = 6'h1d == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_29_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12958 = 6'h1e == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_30_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12959 = 6'h1f == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_31_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12960 = 6'h20 == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_32_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12961 = 6'h21 == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_33_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12962 = 6'h22 == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_34_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12963 = 6'h23 == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_35_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12964 = 6'h24 == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_36_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12965 = 6'h25 == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_37_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12966 = 6'h26 == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_38_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12967 = 6'h27 == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_39_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12968 = 6'h28 == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_40_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12969 = 6'h29 == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_41_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12970 = 6'h2a == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_42_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12971 = 6'h2b == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_43_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12972 = 6'h2c == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_44_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12973 = 6'h2d == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_45_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12974 = 6'h2e == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_46_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12975 = 6'h2f == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_47_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12976 = 6'h30 == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_48_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12977 = 6'h31 == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_49_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12978 = 6'h32 == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_50_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12979 = 6'h33 == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_51_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12980 = 6'h34 == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_52_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12981 = 6'h35 == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_53_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12982 = 6'h36 == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_54_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12983 = 6'h37 == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_55_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12984 = 6'h38 == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_56_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12985 = 6'h39 == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_57_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12986 = 6'h3a == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_58_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12987 = 6'h3b == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_59_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12988 = 6'h3c == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_60_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12989 = 6'h3d == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_61_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12990 = 6'h3e == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_62_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12991 = 6'h3f == allocate_ptr[5:0] ? _rob_uop_T_pc : rob_uop_63_pc; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12992 = 6'h0 == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_0_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12993 = 6'h1 == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_1_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12994 = 6'h2 == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_2_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12995 = 6'h3 == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_3_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12996 = 6'h4 == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_4_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12997 = 6'h5 == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_5_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12998 = 6'h6 == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_6_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_12999 = 6'h7 == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_7_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13000 = 6'h8 == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_8_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13001 = 6'h9 == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_9_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13002 = 6'ha == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_10_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13003 = 6'hb == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_11_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13004 = 6'hc == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_12_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13005 = 6'hd == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_13_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13006 = 6'he == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_14_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13007 = 6'hf == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_15_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13008 = 6'h10 == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_16_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13009 = 6'h11 == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_17_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13010 = 6'h12 == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_18_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13011 = 6'h13 == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_19_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13012 = 6'h14 == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_20_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13013 = 6'h15 == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_21_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13014 = 6'h16 == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_22_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13015 = 6'h17 == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_23_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13016 = 6'h18 == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_24_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13017 = 6'h19 == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_25_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13018 = 6'h1a == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_26_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13019 = 6'h1b == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_27_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13020 = 6'h1c == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_28_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13021 = 6'h1d == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_29_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13022 = 6'h1e == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_30_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13023 = 6'h1f == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_31_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13024 = 6'h20 == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_32_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13025 = 6'h21 == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_33_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13026 = 6'h22 == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_34_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13027 = 6'h23 == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_35_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13028 = 6'h24 == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_36_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13029 = 6'h25 == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_37_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13030 = 6'h26 == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_38_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13031 = 6'h27 == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_39_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13032 = 6'h28 == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_40_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13033 = 6'h29 == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_41_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13034 = 6'h2a == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_42_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13035 = 6'h2b == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_43_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13036 = 6'h2c == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_44_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13037 = 6'h2d == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_45_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13038 = 6'h2e == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_46_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13039 = 6'h2f == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_47_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13040 = 6'h30 == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_48_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13041 = 6'h31 == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_49_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13042 = 6'h32 == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_50_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13043 = 6'h33 == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_51_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13044 = 6'h34 == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_52_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13045 = 6'h35 == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_53_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13046 = 6'h36 == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_54_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13047 = 6'h37 == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_55_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13048 = 6'h38 == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_56_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13049 = 6'h39 == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_57_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13050 = 6'h3a == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_58_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13051 = 6'h3b == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_59_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13052 = 6'h3c == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_60_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13053 = 6'h3d == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_61_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13054 = 6'h3e == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_62_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_13055 = 6'h3f == allocate_ptr[5:0] ? _rob_uop_T_inst : rob_uop_63_inst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13056 = 6'h0 == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_0_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13057 = 6'h1 == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_1_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13058 = 6'h2 == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_2_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13059 = 6'h3 == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_3_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13060 = 6'h4 == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_4_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13061 = 6'h5 == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_5_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13062 = 6'h6 == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_6_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13063 = 6'h7 == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_7_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13064 = 6'h8 == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_8_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13065 = 6'h9 == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_9_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13066 = 6'ha == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_10_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13067 = 6'hb == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_11_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13068 = 6'hc == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_12_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13069 = 6'hd == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_13_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13070 = 6'he == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_14_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13071 = 6'hf == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_15_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13072 = 6'h10 == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_16_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13073 = 6'h11 == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_17_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13074 = 6'h12 == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_18_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13075 = 6'h13 == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_19_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13076 = 6'h14 == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_20_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13077 = 6'h15 == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_21_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13078 = 6'h16 == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_22_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13079 = 6'h17 == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_23_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13080 = 6'h18 == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_24_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13081 = 6'h19 == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_25_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13082 = 6'h1a == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_26_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13083 = 6'h1b == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_27_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13084 = 6'h1c == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_28_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13085 = 6'h1d == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_29_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13086 = 6'h1e == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_30_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13087 = 6'h1f == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_31_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13088 = 6'h20 == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_32_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13089 = 6'h21 == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_33_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13090 = 6'h22 == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_34_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13091 = 6'h23 == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_35_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13092 = 6'h24 == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_36_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13093 = 6'h25 == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_37_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13094 = 6'h26 == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_38_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13095 = 6'h27 == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_39_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13096 = 6'h28 == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_40_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13097 = 6'h29 == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_41_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13098 = 6'h2a == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_42_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13099 = 6'h2b == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_43_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13100 = 6'h2c == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_44_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13101 = 6'h2d == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_45_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13102 = 6'h2e == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_46_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13103 = 6'h2f == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_47_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13104 = 6'h30 == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_48_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13105 = 6'h31 == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_49_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13106 = 6'h32 == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_50_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13107 = 6'h33 == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_51_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13108 = 6'h34 == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_52_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13109 = 6'h35 == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_53_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13110 = 6'h36 == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_54_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13111 = 6'h37 == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_55_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13112 = 6'h38 == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_56_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13113 = 6'h39 == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_57_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13114 = 6'h3a == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_58_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13115 = 6'h3b == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_59_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13116 = 6'h3c == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_60_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13117 = 6'h3d == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_61_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13118 = 6'h3e == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_62_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13119 = 6'h3f == allocate_ptr[5:0] ? _rob_uop_T_func_code : rob_uop_63_func_code; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13440 = 6'h0 == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_0_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13441 = 6'h1 == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_1_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13442 = 6'h2 == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_2_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13443 = 6'h3 == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_3_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13444 = 6'h4 == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_4_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13445 = 6'h5 == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_5_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13446 = 6'h6 == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_6_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13447 = 6'h7 == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_7_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13448 = 6'h8 == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_8_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13449 = 6'h9 == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_9_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13450 = 6'ha == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_10_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13451 = 6'hb == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_11_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13452 = 6'hc == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_12_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13453 = 6'hd == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_13_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13454 = 6'he == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_14_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13455 = 6'hf == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_15_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13456 = 6'h10 == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_16_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13457 = 6'h11 == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_17_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13458 = 6'h12 == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_18_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13459 = 6'h13 == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_19_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13460 = 6'h14 == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_20_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13461 = 6'h15 == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_21_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13462 = 6'h16 == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_22_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13463 = 6'h17 == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_23_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13464 = 6'h18 == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_24_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13465 = 6'h19 == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_25_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13466 = 6'h1a == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_26_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13467 = 6'h1b == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_27_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13468 = 6'h1c == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_28_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13469 = 6'h1d == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_29_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13470 = 6'h1e == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_30_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13471 = 6'h1f == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_31_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13472 = 6'h20 == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_32_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13473 = 6'h21 == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_33_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13474 = 6'h22 == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_34_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13475 = 6'h23 == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_35_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13476 = 6'h24 == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_36_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13477 = 6'h25 == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_37_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13478 = 6'h26 == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_38_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13479 = 6'h27 == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_39_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13480 = 6'h28 == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_40_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13481 = 6'h29 == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_41_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13482 = 6'h2a == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_42_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13483 = 6'h2b == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_43_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13484 = 6'h2c == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_44_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13485 = 6'h2d == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_45_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13486 = 6'h2e == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_46_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13487 = 6'h2f == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_47_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13488 = 6'h30 == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_48_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13489 = 6'h31 == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_49_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13490 = 6'h32 == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_50_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13491 = 6'h33 == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_51_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13492 = 6'h34 == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_52_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13493 = 6'h35 == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_53_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13494 = 6'h36 == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_54_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13495 = 6'h37 == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_55_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13496 = 6'h38 == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_56_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13497 = 6'h39 == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_57_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13498 = 6'h3a == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_58_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13499 = 6'h3b == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_59_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13500 = 6'h3c == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_60_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13501 = 6'h3d == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_61_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13502 = 6'h3e == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_62_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13503 = 6'h3f == allocate_ptr[5:0] ? _rob_uop_T_phy_dst : rob_uop_63_phy_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13504 = 6'h0 == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_0_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13505 = 6'h1 == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_1_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13506 = 6'h2 == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_2_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13507 = 6'h3 == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_3_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13508 = 6'h4 == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_4_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13509 = 6'h5 == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_5_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13510 = 6'h6 == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_6_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13511 = 6'h7 == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_7_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13512 = 6'h8 == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_8_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13513 = 6'h9 == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_9_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13514 = 6'ha == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_10_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13515 = 6'hb == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_11_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13516 = 6'hc == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_12_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13517 = 6'hd == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_13_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13518 = 6'he == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_14_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13519 = 6'hf == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_15_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13520 = 6'h10 == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_16_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13521 = 6'h11 == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_17_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13522 = 6'h12 == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_18_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13523 = 6'h13 == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_19_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13524 = 6'h14 == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_20_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13525 = 6'h15 == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_21_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13526 = 6'h16 == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_22_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13527 = 6'h17 == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_23_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13528 = 6'h18 == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_24_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13529 = 6'h19 == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_25_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13530 = 6'h1a == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_26_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13531 = 6'h1b == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_27_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13532 = 6'h1c == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_28_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13533 = 6'h1d == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_29_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13534 = 6'h1e == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_30_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13535 = 6'h1f == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_31_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13536 = 6'h20 == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_32_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13537 = 6'h21 == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_33_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13538 = 6'h22 == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_34_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13539 = 6'h23 == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_35_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13540 = 6'h24 == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_36_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13541 = 6'h25 == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_37_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13542 = 6'h26 == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_38_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13543 = 6'h27 == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_39_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13544 = 6'h28 == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_40_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13545 = 6'h29 == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_41_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13546 = 6'h2a == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_42_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13547 = 6'h2b == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_43_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13548 = 6'h2c == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_44_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13549 = 6'h2d == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_45_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13550 = 6'h2e == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_46_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13551 = 6'h2f == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_47_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13552 = 6'h30 == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_48_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13553 = 6'h31 == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_49_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13554 = 6'h32 == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_50_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13555 = 6'h33 == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_51_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13556 = 6'h34 == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_52_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13557 = 6'h35 == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_53_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13558 = 6'h36 == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_54_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13559 = 6'h37 == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_55_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13560 = 6'h38 == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_56_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13561 = 6'h39 == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_57_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13562 = 6'h3a == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_58_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13563 = 6'h3b == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_59_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13564 = 6'h3c == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_60_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13565 = 6'h3d == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_61_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13566 = 6'h3e == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_62_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [6:0] _GEN_13567 = 6'h3f == allocate_ptr[5:0] ? _rob_uop_T_stale_dst : rob_uop_63_stale_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13568 = 6'h0 == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_0_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13569 = 6'h1 == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_1_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13570 = 6'h2 == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_2_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13571 = 6'h3 == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_3_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13572 = 6'h4 == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_4_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13573 = 6'h5 == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_5_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13574 = 6'h6 == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_6_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13575 = 6'h7 == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_7_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13576 = 6'h8 == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_8_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13577 = 6'h9 == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_9_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13578 = 6'ha == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_10_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13579 = 6'hb == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_11_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13580 = 6'hc == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_12_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13581 = 6'hd == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_13_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13582 = 6'he == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_14_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13583 = 6'hf == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_15_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13584 = 6'h10 == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_16_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13585 = 6'h11 == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_17_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13586 = 6'h12 == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_18_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13587 = 6'h13 == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_19_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13588 = 6'h14 == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_20_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13589 = 6'h15 == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_21_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13590 = 6'h16 == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_22_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13591 = 6'h17 == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_23_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13592 = 6'h18 == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_24_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13593 = 6'h19 == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_25_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13594 = 6'h1a == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_26_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13595 = 6'h1b == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_27_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13596 = 6'h1c == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_28_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13597 = 6'h1d == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_29_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13598 = 6'h1e == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_30_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13599 = 6'h1f == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_31_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13600 = 6'h20 == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_32_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13601 = 6'h21 == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_33_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13602 = 6'h22 == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_34_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13603 = 6'h23 == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_35_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13604 = 6'h24 == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_36_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13605 = 6'h25 == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_37_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13606 = 6'h26 == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_38_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13607 = 6'h27 == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_39_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13608 = 6'h28 == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_40_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13609 = 6'h29 == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_41_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13610 = 6'h2a == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_42_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13611 = 6'h2b == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_43_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13612 = 6'h2c == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_44_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13613 = 6'h2d == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_45_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13614 = 6'h2e == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_46_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13615 = 6'h2f == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_47_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13616 = 6'h30 == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_48_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13617 = 6'h31 == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_49_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13618 = 6'h32 == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_50_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13619 = 6'h33 == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_51_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13620 = 6'h34 == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_52_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13621 = 6'h35 == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_53_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13622 = 6'h36 == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_54_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13623 = 6'h37 == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_55_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13624 = 6'h38 == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_56_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13625 = 6'h39 == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_57_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13626 = 6'h3a == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_58_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13627 = 6'h3b == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_59_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13628 = 6'h3c == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_60_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13629 = 6'h3d == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_61_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13630 = 6'h3e == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_62_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_13631 = 6'h3f == allocate_ptr[5:0] ? _rob_uop_T_arch_dst : rob_uop_63_arch_dst; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14336 = 6'h0 == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_0_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14337 = 6'h1 == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_1_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14338 = 6'h2 == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_2_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14339 = 6'h3 == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_3_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14340 = 6'h4 == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_4_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14341 = 6'h5 == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_5_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14342 = 6'h6 == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_6_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14343 = 6'h7 == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_7_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14344 = 6'h8 == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_8_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14345 = 6'h9 == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_9_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14346 = 6'ha == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_10_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14347 = 6'hb == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_11_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14348 = 6'hc == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_12_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14349 = 6'hd == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_13_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14350 = 6'he == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_14_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14351 = 6'hf == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_15_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14352 = 6'h10 == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_16_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14353 = 6'h11 == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_17_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14354 = 6'h12 == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_18_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14355 = 6'h13 == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_19_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14356 = 6'h14 == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_20_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14357 = 6'h15 == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_21_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14358 = 6'h16 == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_22_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14359 = 6'h17 == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_23_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14360 = 6'h18 == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_24_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14361 = 6'h19 == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_25_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14362 = 6'h1a == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_26_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14363 = 6'h1b == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_27_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14364 = 6'h1c == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_28_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14365 = 6'h1d == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_29_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14366 = 6'h1e == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_30_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14367 = 6'h1f == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_31_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14368 = 6'h20 == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_32_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14369 = 6'h21 == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_33_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14370 = 6'h22 == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_34_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14371 = 6'h23 == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_35_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14372 = 6'h24 == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_36_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14373 = 6'h25 == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_37_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14374 = 6'h26 == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_38_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14375 = 6'h27 == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_39_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14376 = 6'h28 == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_40_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14377 = 6'h29 == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_41_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14378 = 6'h2a == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_42_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14379 = 6'h2b == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_43_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14380 = 6'h2c == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_44_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14381 = 6'h2d == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_45_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14382 = 6'h2e == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_46_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14383 = 6'h2f == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_47_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14384 = 6'h30 == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_48_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14385 = 6'h31 == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_49_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14386 = 6'h32 == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_50_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14387 = 6'h33 == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_51_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14388 = 6'h34 == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_52_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14389 = 6'h35 == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_53_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14390 = 6'h36 == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_54_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14391 = 6'h37 == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_55_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14392 = 6'h38 == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_56_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14393 = 6'h39 == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_57_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14394 = 6'h3a == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_58_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14395 = 6'h3b == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_59_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14396 = 6'h3c == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_60_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14397 = 6'h3d == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_61_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14398 = 6'h3e == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_62_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [63:0] _GEN_14399 = 6'h3f == allocate_ptr[5:0] ? _rob_uop_T_src1_value : rob_uop_63_src1_value; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14656 = 6'h0 == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_0_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14657 = 6'h1 == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_1_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14658 = 6'h2 == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_2_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14659 = 6'h3 == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_3_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14660 = 6'h4 == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_4_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14661 = 6'h5 == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_5_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14662 = 6'h6 == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_6_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14663 = 6'h7 == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_7_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14664 = 6'h8 == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_8_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14665 = 6'h9 == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_9_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14666 = 6'ha == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_10_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14667 = 6'hb == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_11_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14668 = 6'hc == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_12_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14669 = 6'hd == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_13_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14670 = 6'he == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_14_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14671 = 6'hf == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_15_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14672 = 6'h10 == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_16_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14673 = 6'h11 == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_17_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14674 = 6'h12 == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_18_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14675 = 6'h13 == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_19_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14676 = 6'h14 == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_20_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14677 = 6'h15 == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_21_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14678 = 6'h16 == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_22_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14679 = 6'h17 == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_23_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14680 = 6'h18 == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_24_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14681 = 6'h19 == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_25_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14682 = 6'h1a == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_26_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14683 = 6'h1b == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_27_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14684 = 6'h1c == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_28_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14685 = 6'h1d == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_29_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14686 = 6'h1e == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_30_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14687 = 6'h1f == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_31_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14688 = 6'h20 == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_32_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14689 = 6'h21 == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_33_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14690 = 6'h22 == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_34_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14691 = 6'h23 == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_35_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14692 = 6'h24 == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_36_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14693 = 6'h25 == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_37_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14694 = 6'h26 == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_38_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14695 = 6'h27 == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_39_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14696 = 6'h28 == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_40_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14697 = 6'h29 == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_41_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14698 = 6'h2a == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_42_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14699 = 6'h2b == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_43_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14700 = 6'h2c == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_44_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14701 = 6'h2d == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_45_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14702 = 6'h2e == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_46_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14703 = 6'h2f == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_47_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14704 = 6'h30 == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_48_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14705 = 6'h31 == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_49_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14706 = 6'h32 == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_50_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14707 = 6'h33 == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_51_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14708 = 6'h34 == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_52_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14709 = 6'h35 == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_53_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14710 = 6'h36 == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_54_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14711 = 6'h37 == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_55_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14712 = 6'h38 == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_56_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14713 = 6'h39 == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_57_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14714 = 6'h3a == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_58_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14715 = 6'h3b == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_59_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14716 = 6'h3c == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_60_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14717 = 6'h3d == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_61_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14718 = 6'h3e == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_62_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [4:0] _GEN_14719 = 6'h3f == allocate_ptr[5:0] ? _rob_uop_T_alu_sel : rob_uop_63_alu_sel; // @[rob.scala 134:{31,31} 82:26]
  wire [31:0] _GEN_15040 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12928 :
    rob_uop_0_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15041 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12929 :
    rob_uop_1_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15042 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12930 :
    rob_uop_2_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15043 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12931 :
    rob_uop_3_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15044 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12932 :
    rob_uop_4_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15045 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12933 :
    rob_uop_5_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15046 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12934 :
    rob_uop_6_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15047 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12935 :
    rob_uop_7_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15048 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12936 :
    rob_uop_8_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15049 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12937 :
    rob_uop_9_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15050 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12938 :
    rob_uop_10_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15051 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12939 :
    rob_uop_11_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15052 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12940 :
    rob_uop_12_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15053 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12941 :
    rob_uop_13_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15054 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12942 :
    rob_uop_14_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15055 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12943 :
    rob_uop_15_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15056 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12944 :
    rob_uop_16_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15057 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12945 :
    rob_uop_17_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15058 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12946 :
    rob_uop_18_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15059 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12947 :
    rob_uop_19_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15060 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12948 :
    rob_uop_20_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15061 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12949 :
    rob_uop_21_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15062 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12950 :
    rob_uop_22_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15063 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12951 :
    rob_uop_23_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15064 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12952 :
    rob_uop_24_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15065 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12953 :
    rob_uop_25_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15066 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12954 :
    rob_uop_26_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15067 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12955 :
    rob_uop_27_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15068 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12956 :
    rob_uop_28_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15069 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12957 :
    rob_uop_29_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15070 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12958 :
    rob_uop_30_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15071 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12959 :
    rob_uop_31_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15072 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12960 :
    rob_uop_32_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15073 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12961 :
    rob_uop_33_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15074 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12962 :
    rob_uop_34_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15075 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12963 :
    rob_uop_35_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15076 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12964 :
    rob_uop_36_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15077 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12965 :
    rob_uop_37_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15078 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12966 :
    rob_uop_38_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15079 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12967 :
    rob_uop_39_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15080 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12968 :
    rob_uop_40_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15081 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12969 :
    rob_uop_41_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15082 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12970 :
    rob_uop_42_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15083 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12971 :
    rob_uop_43_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15084 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12972 :
    rob_uop_44_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15085 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12973 :
    rob_uop_45_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15086 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12974 :
    rob_uop_46_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15087 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12975 :
    rob_uop_47_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15088 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12976 :
    rob_uop_48_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15089 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12977 :
    rob_uop_49_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15090 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12978 :
    rob_uop_50_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15091 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12979 :
    rob_uop_51_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15092 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12980 :
    rob_uop_52_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15093 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12981 :
    rob_uop_53_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15094 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12982 :
    rob_uop_54_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15095 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12983 :
    rob_uop_55_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15096 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12984 :
    rob_uop_56_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15097 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12985 :
    rob_uop_57_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15098 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12986 :
    rob_uop_58_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15099 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12987 :
    rob_uop_59_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15100 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12988 :
    rob_uop_60_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15101 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12989 :
    rob_uop_61_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15102 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12990 :
    rob_uop_62_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15103 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12991 :
    rob_uop_63_pc; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15104 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12992 :
    rob_uop_0_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15105 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12993 :
    rob_uop_1_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15106 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12994 :
    rob_uop_2_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15107 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12995 :
    rob_uop_3_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15108 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12996 :
    rob_uop_4_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15109 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12997 :
    rob_uop_5_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15110 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12998 :
    rob_uop_6_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15111 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_12999 :
    rob_uop_7_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15112 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13000 :
    rob_uop_8_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15113 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13001 :
    rob_uop_9_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15114 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13002 :
    rob_uop_10_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15115 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13003 :
    rob_uop_11_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15116 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13004 :
    rob_uop_12_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15117 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13005 :
    rob_uop_13_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15118 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13006 :
    rob_uop_14_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15119 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13007 :
    rob_uop_15_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15120 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13008 :
    rob_uop_16_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15121 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13009 :
    rob_uop_17_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15122 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13010 :
    rob_uop_18_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15123 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13011 :
    rob_uop_19_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15124 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13012 :
    rob_uop_20_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15125 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13013 :
    rob_uop_21_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15126 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13014 :
    rob_uop_22_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15127 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13015 :
    rob_uop_23_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15128 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13016 :
    rob_uop_24_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15129 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13017 :
    rob_uop_25_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15130 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13018 :
    rob_uop_26_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15131 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13019 :
    rob_uop_27_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15132 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13020 :
    rob_uop_28_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15133 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13021 :
    rob_uop_29_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15134 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13022 :
    rob_uop_30_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15135 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13023 :
    rob_uop_31_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15136 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13024 :
    rob_uop_32_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15137 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13025 :
    rob_uop_33_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15138 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13026 :
    rob_uop_34_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15139 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13027 :
    rob_uop_35_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15140 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13028 :
    rob_uop_36_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15141 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13029 :
    rob_uop_37_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15142 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13030 :
    rob_uop_38_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15143 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13031 :
    rob_uop_39_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15144 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13032 :
    rob_uop_40_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15145 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13033 :
    rob_uop_41_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15146 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13034 :
    rob_uop_42_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15147 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13035 :
    rob_uop_43_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15148 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13036 :
    rob_uop_44_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15149 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13037 :
    rob_uop_45_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15150 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13038 :
    rob_uop_46_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15151 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13039 :
    rob_uop_47_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15152 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13040 :
    rob_uop_48_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15153 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13041 :
    rob_uop_49_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15154 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13042 :
    rob_uop_50_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15155 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13043 :
    rob_uop_51_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15156 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13044 :
    rob_uop_52_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15157 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13045 :
    rob_uop_53_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15158 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13046 :
    rob_uop_54_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15159 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13047 :
    rob_uop_55_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15160 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13048 :
    rob_uop_56_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15161 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13049 :
    rob_uop_57_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15162 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13050 :
    rob_uop_58_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15163 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13051 :
    rob_uop_59_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15164 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13052 :
    rob_uop_60_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15165 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13053 :
    rob_uop_61_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15166 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13054 :
    rob_uop_62_inst; // @[rob.scala 133:89 82:26]
  wire [31:0] _GEN_15167 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13055 :
    rob_uop_63_inst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15168 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13056 :
    rob_uop_0_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15169 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13057 :
    rob_uop_1_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15170 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13058 :
    rob_uop_2_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15171 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13059 :
    rob_uop_3_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15172 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13060 :
    rob_uop_4_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15173 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13061 :
    rob_uop_5_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15174 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13062 :
    rob_uop_6_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15175 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13063 :
    rob_uop_7_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15176 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13064 :
    rob_uop_8_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15177 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13065 :
    rob_uop_9_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15178 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13066 :
    rob_uop_10_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15179 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13067 :
    rob_uop_11_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15180 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13068 :
    rob_uop_12_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15181 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13069 :
    rob_uop_13_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15182 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13070 :
    rob_uop_14_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15183 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13071 :
    rob_uop_15_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15184 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13072 :
    rob_uop_16_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15185 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13073 :
    rob_uop_17_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15186 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13074 :
    rob_uop_18_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15187 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13075 :
    rob_uop_19_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15188 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13076 :
    rob_uop_20_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15189 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13077 :
    rob_uop_21_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15190 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13078 :
    rob_uop_22_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15191 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13079 :
    rob_uop_23_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15192 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13080 :
    rob_uop_24_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15193 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13081 :
    rob_uop_25_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15194 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13082 :
    rob_uop_26_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15195 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13083 :
    rob_uop_27_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15196 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13084 :
    rob_uop_28_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15197 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13085 :
    rob_uop_29_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15198 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13086 :
    rob_uop_30_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15199 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13087 :
    rob_uop_31_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15200 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13088 :
    rob_uop_32_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15201 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13089 :
    rob_uop_33_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15202 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13090 :
    rob_uop_34_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15203 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13091 :
    rob_uop_35_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15204 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13092 :
    rob_uop_36_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15205 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13093 :
    rob_uop_37_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15206 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13094 :
    rob_uop_38_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15207 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13095 :
    rob_uop_39_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15208 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13096 :
    rob_uop_40_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15209 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13097 :
    rob_uop_41_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15210 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13098 :
    rob_uop_42_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15211 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13099 :
    rob_uop_43_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15212 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13100 :
    rob_uop_44_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15213 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13101 :
    rob_uop_45_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15214 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13102 :
    rob_uop_46_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15215 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13103 :
    rob_uop_47_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15216 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13104 :
    rob_uop_48_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15217 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13105 :
    rob_uop_49_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15218 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13106 :
    rob_uop_50_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15219 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13107 :
    rob_uop_51_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15220 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13108 :
    rob_uop_52_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15221 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13109 :
    rob_uop_53_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15222 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13110 :
    rob_uop_54_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15223 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13111 :
    rob_uop_55_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15224 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13112 :
    rob_uop_56_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15225 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13113 :
    rob_uop_57_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15226 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13114 :
    rob_uop_58_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15227 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13115 :
    rob_uop_59_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15228 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13116 :
    rob_uop_60_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15229 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13117 :
    rob_uop_61_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15230 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13118 :
    rob_uop_62_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15231 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13119 :
    rob_uop_63_func_code; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15552 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13440 :
    rob_uop_0_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15553 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13441 :
    rob_uop_1_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15554 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13442 :
    rob_uop_2_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15555 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13443 :
    rob_uop_3_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15556 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13444 :
    rob_uop_4_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15557 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13445 :
    rob_uop_5_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15558 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13446 :
    rob_uop_6_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15559 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13447 :
    rob_uop_7_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15560 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13448 :
    rob_uop_8_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15561 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13449 :
    rob_uop_9_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15562 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13450 :
    rob_uop_10_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15563 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13451 :
    rob_uop_11_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15564 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13452 :
    rob_uop_12_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15565 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13453 :
    rob_uop_13_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15566 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13454 :
    rob_uop_14_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15567 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13455 :
    rob_uop_15_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15568 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13456 :
    rob_uop_16_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15569 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13457 :
    rob_uop_17_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15570 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13458 :
    rob_uop_18_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15571 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13459 :
    rob_uop_19_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15572 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13460 :
    rob_uop_20_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15573 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13461 :
    rob_uop_21_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15574 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13462 :
    rob_uop_22_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15575 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13463 :
    rob_uop_23_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15576 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13464 :
    rob_uop_24_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15577 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13465 :
    rob_uop_25_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15578 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13466 :
    rob_uop_26_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15579 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13467 :
    rob_uop_27_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15580 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13468 :
    rob_uop_28_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15581 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13469 :
    rob_uop_29_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15582 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13470 :
    rob_uop_30_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15583 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13471 :
    rob_uop_31_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15584 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13472 :
    rob_uop_32_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15585 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13473 :
    rob_uop_33_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15586 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13474 :
    rob_uop_34_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15587 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13475 :
    rob_uop_35_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15588 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13476 :
    rob_uop_36_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15589 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13477 :
    rob_uop_37_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15590 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13478 :
    rob_uop_38_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15591 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13479 :
    rob_uop_39_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15592 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13480 :
    rob_uop_40_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15593 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13481 :
    rob_uop_41_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15594 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13482 :
    rob_uop_42_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15595 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13483 :
    rob_uop_43_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15596 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13484 :
    rob_uop_44_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15597 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13485 :
    rob_uop_45_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15598 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13486 :
    rob_uop_46_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15599 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13487 :
    rob_uop_47_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15600 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13488 :
    rob_uop_48_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15601 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13489 :
    rob_uop_49_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15602 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13490 :
    rob_uop_50_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15603 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13491 :
    rob_uop_51_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15604 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13492 :
    rob_uop_52_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15605 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13493 :
    rob_uop_53_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15606 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13494 :
    rob_uop_54_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15607 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13495 :
    rob_uop_55_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15608 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13496 :
    rob_uop_56_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15609 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13497 :
    rob_uop_57_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15610 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13498 :
    rob_uop_58_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15611 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13499 :
    rob_uop_59_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15612 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13500 :
    rob_uop_60_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15613 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13501 :
    rob_uop_61_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15614 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13502 :
    rob_uop_62_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15615 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13503 :
    rob_uop_63_phy_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15616 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13504 :
    rob_uop_0_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15617 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13505 :
    rob_uop_1_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15618 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13506 :
    rob_uop_2_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15619 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13507 :
    rob_uop_3_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15620 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13508 :
    rob_uop_4_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15621 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13509 :
    rob_uop_5_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15622 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13510 :
    rob_uop_6_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15623 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13511 :
    rob_uop_7_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15624 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13512 :
    rob_uop_8_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15625 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13513 :
    rob_uop_9_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15626 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13514 :
    rob_uop_10_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15627 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13515 :
    rob_uop_11_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15628 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13516 :
    rob_uop_12_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15629 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13517 :
    rob_uop_13_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15630 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13518 :
    rob_uop_14_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15631 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13519 :
    rob_uop_15_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15632 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13520 :
    rob_uop_16_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15633 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13521 :
    rob_uop_17_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15634 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13522 :
    rob_uop_18_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15635 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13523 :
    rob_uop_19_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15636 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13524 :
    rob_uop_20_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15637 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13525 :
    rob_uop_21_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15638 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13526 :
    rob_uop_22_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15639 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13527 :
    rob_uop_23_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15640 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13528 :
    rob_uop_24_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15641 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13529 :
    rob_uop_25_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15642 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13530 :
    rob_uop_26_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15643 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13531 :
    rob_uop_27_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15644 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13532 :
    rob_uop_28_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15645 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13533 :
    rob_uop_29_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15646 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13534 :
    rob_uop_30_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15647 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13535 :
    rob_uop_31_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15648 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13536 :
    rob_uop_32_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15649 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13537 :
    rob_uop_33_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15650 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13538 :
    rob_uop_34_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15651 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13539 :
    rob_uop_35_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15652 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13540 :
    rob_uop_36_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15653 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13541 :
    rob_uop_37_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15654 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13542 :
    rob_uop_38_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15655 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13543 :
    rob_uop_39_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15656 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13544 :
    rob_uop_40_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15657 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13545 :
    rob_uop_41_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15658 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13546 :
    rob_uop_42_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15659 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13547 :
    rob_uop_43_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15660 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13548 :
    rob_uop_44_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15661 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13549 :
    rob_uop_45_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15662 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13550 :
    rob_uop_46_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15663 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13551 :
    rob_uop_47_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15664 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13552 :
    rob_uop_48_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15665 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13553 :
    rob_uop_49_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15666 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13554 :
    rob_uop_50_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15667 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13555 :
    rob_uop_51_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15668 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13556 :
    rob_uop_52_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15669 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13557 :
    rob_uop_53_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15670 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13558 :
    rob_uop_54_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15671 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13559 :
    rob_uop_55_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15672 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13560 :
    rob_uop_56_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15673 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13561 :
    rob_uop_57_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15674 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13562 :
    rob_uop_58_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15675 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13563 :
    rob_uop_59_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15676 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13564 :
    rob_uop_60_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15677 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13565 :
    rob_uop_61_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15678 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13566 :
    rob_uop_62_stale_dst; // @[rob.scala 133:89 82:26]
  wire [6:0] _GEN_15679 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13567 :
    rob_uop_63_stale_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15680 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13568 :
    rob_uop_0_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15681 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13569 :
    rob_uop_1_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15682 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13570 :
    rob_uop_2_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15683 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13571 :
    rob_uop_3_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15684 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13572 :
    rob_uop_4_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15685 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13573 :
    rob_uop_5_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15686 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13574 :
    rob_uop_6_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15687 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13575 :
    rob_uop_7_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15688 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13576 :
    rob_uop_8_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15689 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13577 :
    rob_uop_9_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15690 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13578 :
    rob_uop_10_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15691 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13579 :
    rob_uop_11_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15692 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13580 :
    rob_uop_12_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15693 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13581 :
    rob_uop_13_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15694 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13582 :
    rob_uop_14_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15695 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13583 :
    rob_uop_15_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15696 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13584 :
    rob_uop_16_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15697 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13585 :
    rob_uop_17_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15698 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13586 :
    rob_uop_18_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15699 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13587 :
    rob_uop_19_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15700 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13588 :
    rob_uop_20_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15701 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13589 :
    rob_uop_21_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15702 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13590 :
    rob_uop_22_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15703 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13591 :
    rob_uop_23_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15704 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13592 :
    rob_uop_24_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15705 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13593 :
    rob_uop_25_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15706 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13594 :
    rob_uop_26_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15707 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13595 :
    rob_uop_27_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15708 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13596 :
    rob_uop_28_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15709 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13597 :
    rob_uop_29_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15710 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13598 :
    rob_uop_30_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15711 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13599 :
    rob_uop_31_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15712 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13600 :
    rob_uop_32_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15713 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13601 :
    rob_uop_33_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15714 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13602 :
    rob_uop_34_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15715 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13603 :
    rob_uop_35_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15716 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13604 :
    rob_uop_36_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15717 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13605 :
    rob_uop_37_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15718 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13606 :
    rob_uop_38_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15719 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13607 :
    rob_uop_39_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15720 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13608 :
    rob_uop_40_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15721 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13609 :
    rob_uop_41_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15722 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13610 :
    rob_uop_42_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15723 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13611 :
    rob_uop_43_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15724 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13612 :
    rob_uop_44_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15725 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13613 :
    rob_uop_45_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15726 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13614 :
    rob_uop_46_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15727 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13615 :
    rob_uop_47_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15728 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13616 :
    rob_uop_48_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15729 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13617 :
    rob_uop_49_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15730 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13618 :
    rob_uop_50_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15731 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13619 :
    rob_uop_51_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15732 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13620 :
    rob_uop_52_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15733 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13621 :
    rob_uop_53_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15734 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13622 :
    rob_uop_54_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15735 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13623 :
    rob_uop_55_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15736 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13624 :
    rob_uop_56_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15737 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13625 :
    rob_uop_57_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15738 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13626 :
    rob_uop_58_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15739 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13627 :
    rob_uop_59_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15740 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13628 :
    rob_uop_60_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15741 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13629 :
    rob_uop_61_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15742 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13630 :
    rob_uop_62_arch_dst; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_15743 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_13631 :
    rob_uop_63_arch_dst; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16384 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10048 :
    rob_uop_0_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16385 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10049 :
    rob_uop_1_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16386 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10050 :
    rob_uop_2_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16387 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10051 :
    rob_uop_3_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16388 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10052 :
    rob_uop_4_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16389 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10053 :
    rob_uop_5_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16390 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10054 :
    rob_uop_6_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16391 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10055 :
    rob_uop_7_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16392 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10056 :
    rob_uop_8_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16393 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10057 :
    rob_uop_9_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16394 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10058 :
    rob_uop_10_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16395 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10059 :
    rob_uop_11_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16396 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10060 :
    rob_uop_12_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16397 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10061 :
    rob_uop_13_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16398 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10062 :
    rob_uop_14_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16399 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10063 :
    rob_uop_15_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16400 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10064 :
    rob_uop_16_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16401 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10065 :
    rob_uop_17_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16402 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10066 :
    rob_uop_18_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16403 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10067 :
    rob_uop_19_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16404 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10068 :
    rob_uop_20_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16405 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10069 :
    rob_uop_21_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16406 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10070 :
    rob_uop_22_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16407 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10071 :
    rob_uop_23_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16408 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10072 :
    rob_uop_24_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16409 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10073 :
    rob_uop_25_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16410 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10074 :
    rob_uop_26_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16411 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10075 :
    rob_uop_27_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16412 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10076 :
    rob_uop_28_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16413 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10077 :
    rob_uop_29_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16414 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10078 :
    rob_uop_30_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16415 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10079 :
    rob_uop_31_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16416 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10080 :
    rob_uop_32_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16417 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10081 :
    rob_uop_33_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16418 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10082 :
    rob_uop_34_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16419 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10083 :
    rob_uop_35_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16420 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10084 :
    rob_uop_36_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16421 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10085 :
    rob_uop_37_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16422 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10086 :
    rob_uop_38_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16423 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10087 :
    rob_uop_39_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16424 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10088 :
    rob_uop_40_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16425 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10089 :
    rob_uop_41_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16426 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10090 :
    rob_uop_42_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16427 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10091 :
    rob_uop_43_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16428 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10092 :
    rob_uop_44_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16429 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10093 :
    rob_uop_45_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16430 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10094 :
    rob_uop_46_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16431 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10095 :
    rob_uop_47_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16432 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10096 :
    rob_uop_48_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16433 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10097 :
    rob_uop_49_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16434 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10098 :
    rob_uop_50_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16435 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10099 :
    rob_uop_51_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16436 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10100 :
    rob_uop_52_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16437 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10101 :
    rob_uop_53_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16438 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10102 :
    rob_uop_54_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16439 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10103 :
    rob_uop_55_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16440 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10104 :
    rob_uop_56_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16441 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10105 :
    rob_uop_57_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16442 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10106 :
    rob_uop_58_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16443 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10107 :
    rob_uop_59_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16444 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10108 :
    rob_uop_60_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16445 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10109 :
    rob_uop_61_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16446 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10110 :
    rob_uop_62_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16447 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10111 :
    rob_uop_63_dst_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16448 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14336 :
    rob_uop_0_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16449 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14337 :
    rob_uop_1_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16450 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14338 :
    rob_uop_2_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16451 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14339 :
    rob_uop_3_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16452 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14340 :
    rob_uop_4_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16453 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14341 :
    rob_uop_5_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16454 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14342 :
    rob_uop_6_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16455 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14343 :
    rob_uop_7_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16456 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14344 :
    rob_uop_8_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16457 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14345 :
    rob_uop_9_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16458 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14346 :
    rob_uop_10_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16459 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14347 :
    rob_uop_11_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16460 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14348 :
    rob_uop_12_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16461 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14349 :
    rob_uop_13_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16462 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14350 :
    rob_uop_14_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16463 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14351 :
    rob_uop_15_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16464 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14352 :
    rob_uop_16_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16465 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14353 :
    rob_uop_17_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16466 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14354 :
    rob_uop_18_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16467 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14355 :
    rob_uop_19_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16468 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14356 :
    rob_uop_20_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16469 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14357 :
    rob_uop_21_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16470 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14358 :
    rob_uop_22_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16471 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14359 :
    rob_uop_23_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16472 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14360 :
    rob_uop_24_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16473 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14361 :
    rob_uop_25_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16474 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14362 :
    rob_uop_26_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16475 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14363 :
    rob_uop_27_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16476 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14364 :
    rob_uop_28_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16477 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14365 :
    rob_uop_29_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16478 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14366 :
    rob_uop_30_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16479 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14367 :
    rob_uop_31_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16480 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14368 :
    rob_uop_32_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16481 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14369 :
    rob_uop_33_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16482 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14370 :
    rob_uop_34_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16483 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14371 :
    rob_uop_35_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16484 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14372 :
    rob_uop_36_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16485 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14373 :
    rob_uop_37_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16486 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14374 :
    rob_uop_38_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16487 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14375 :
    rob_uop_39_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16488 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14376 :
    rob_uop_40_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16489 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14377 :
    rob_uop_41_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16490 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14378 :
    rob_uop_42_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16491 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14379 :
    rob_uop_43_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16492 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14380 :
    rob_uop_44_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16493 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14381 :
    rob_uop_45_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16494 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14382 :
    rob_uop_46_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16495 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14383 :
    rob_uop_47_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16496 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14384 :
    rob_uop_48_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16497 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14385 :
    rob_uop_49_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16498 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14386 :
    rob_uop_50_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16499 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14387 :
    rob_uop_51_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16500 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14388 :
    rob_uop_52_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16501 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14389 :
    rob_uop_53_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16502 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14390 :
    rob_uop_54_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16503 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14391 :
    rob_uop_55_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16504 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14392 :
    rob_uop_56_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16505 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14393 :
    rob_uop_57_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16506 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14394 :
    rob_uop_58_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16507 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14395 :
    rob_uop_59_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16508 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14396 :
    rob_uop_60_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16509 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14397 :
    rob_uop_61_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16510 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14398 :
    rob_uop_62_src1_value; // @[rob.scala 133:89 82:26]
  wire [63:0] _GEN_16511 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14399 :
    rob_uop_63_src1_value; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16768 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14656 :
    rob_uop_0_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16769 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14657 :
    rob_uop_1_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16770 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14658 :
    rob_uop_2_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16771 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14659 :
    rob_uop_3_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16772 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14660 :
    rob_uop_4_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16773 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14661 :
    rob_uop_5_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16774 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14662 :
    rob_uop_6_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16775 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14663 :
    rob_uop_7_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16776 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14664 :
    rob_uop_8_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16777 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14665 :
    rob_uop_9_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16778 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14666 :
    rob_uop_10_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16779 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14667 :
    rob_uop_11_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16780 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14668 :
    rob_uop_12_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16781 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14669 :
    rob_uop_13_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16782 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14670 :
    rob_uop_14_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16783 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14671 :
    rob_uop_15_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16784 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14672 :
    rob_uop_16_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16785 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14673 :
    rob_uop_17_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16786 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14674 :
    rob_uop_18_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16787 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14675 :
    rob_uop_19_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16788 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14676 :
    rob_uop_20_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16789 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14677 :
    rob_uop_21_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16790 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14678 :
    rob_uop_22_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16791 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14679 :
    rob_uop_23_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16792 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14680 :
    rob_uop_24_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16793 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14681 :
    rob_uop_25_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16794 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14682 :
    rob_uop_26_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16795 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14683 :
    rob_uop_27_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16796 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14684 :
    rob_uop_28_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16797 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14685 :
    rob_uop_29_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16798 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14686 :
    rob_uop_30_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16799 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14687 :
    rob_uop_31_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16800 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14688 :
    rob_uop_32_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16801 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14689 :
    rob_uop_33_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16802 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14690 :
    rob_uop_34_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16803 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14691 :
    rob_uop_35_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16804 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14692 :
    rob_uop_36_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16805 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14693 :
    rob_uop_37_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16806 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14694 :
    rob_uop_38_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16807 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14695 :
    rob_uop_39_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16808 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14696 :
    rob_uop_40_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16809 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14697 :
    rob_uop_41_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16810 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14698 :
    rob_uop_42_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16811 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14699 :
    rob_uop_43_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16812 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14700 :
    rob_uop_44_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16813 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14701 :
    rob_uop_45_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16814 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14702 :
    rob_uop_46_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16815 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14703 :
    rob_uop_47_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16816 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14704 :
    rob_uop_48_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16817 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14705 :
    rob_uop_49_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16818 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14706 :
    rob_uop_50_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16819 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14707 :
    rob_uop_51_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16820 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14708 :
    rob_uop_52_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16821 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14709 :
    rob_uop_53_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16822 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14710 :
    rob_uop_54_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16823 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14711 :
    rob_uop_55_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16824 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14712 :
    rob_uop_56_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16825 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14713 :
    rob_uop_57_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16826 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14714 :
    rob_uop_58_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16827 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14715 :
    rob_uop_59_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16828 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14716 :
    rob_uop_60_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16829 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14717 :
    rob_uop_61_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16830 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14718 :
    rob_uop_62_alu_sel; // @[rob.scala 133:89 82:26]
  wire [4:0] _GEN_16831 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_14719 :
    rob_uop_63_alu_sel; // @[rob.scala 133:89 82:26]
  wire  _GEN_16960 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10624 : rob_valid_0; // @[rob.scala 133:89 81:28]
  wire  _GEN_16961 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10625 : rob_valid_1; // @[rob.scala 133:89 81:28]
  wire  _GEN_16962 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10626 : rob_valid_2; // @[rob.scala 133:89 81:28]
  wire  _GEN_16963 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10627 : rob_valid_3; // @[rob.scala 133:89 81:28]
  wire  _GEN_16964 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10628 : rob_valid_4; // @[rob.scala 133:89 81:28]
  wire  _GEN_16965 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10629 : rob_valid_5; // @[rob.scala 133:89 81:28]
  wire  _GEN_16966 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10630 : rob_valid_6; // @[rob.scala 133:89 81:28]
  wire  _GEN_16967 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10631 : rob_valid_7; // @[rob.scala 133:89 81:28]
  wire  _GEN_16968 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10632 : rob_valid_8; // @[rob.scala 133:89 81:28]
  wire  _GEN_16969 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10633 : rob_valid_9; // @[rob.scala 133:89 81:28]
  wire  _GEN_16970 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10634 : rob_valid_10; // @[rob.scala 133:89 81:28]
  wire  _GEN_16971 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10635 : rob_valid_11; // @[rob.scala 133:89 81:28]
  wire  _GEN_16972 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10636 : rob_valid_12; // @[rob.scala 133:89 81:28]
  wire  _GEN_16973 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10637 : rob_valid_13; // @[rob.scala 133:89 81:28]
  wire  _GEN_16974 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10638 : rob_valid_14; // @[rob.scala 133:89 81:28]
  wire  _GEN_16975 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10639 : rob_valid_15; // @[rob.scala 133:89 81:28]
  wire  _GEN_16976 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10640 : rob_valid_16; // @[rob.scala 133:89 81:28]
  wire  _GEN_16977 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10641 : rob_valid_17; // @[rob.scala 133:89 81:28]
  wire  _GEN_16978 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10642 : rob_valid_18; // @[rob.scala 133:89 81:28]
  wire  _GEN_16979 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10643 : rob_valid_19; // @[rob.scala 133:89 81:28]
  wire  _GEN_16980 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10644 : rob_valid_20; // @[rob.scala 133:89 81:28]
  wire  _GEN_16981 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10645 : rob_valid_21; // @[rob.scala 133:89 81:28]
  wire  _GEN_16982 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10646 : rob_valid_22; // @[rob.scala 133:89 81:28]
  wire  _GEN_16983 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10647 : rob_valid_23; // @[rob.scala 133:89 81:28]
  wire  _GEN_16984 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10648 : rob_valid_24; // @[rob.scala 133:89 81:28]
  wire  _GEN_16985 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10649 : rob_valid_25; // @[rob.scala 133:89 81:28]
  wire  _GEN_16986 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10650 : rob_valid_26; // @[rob.scala 133:89 81:28]
  wire  _GEN_16987 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10651 : rob_valid_27; // @[rob.scala 133:89 81:28]
  wire  _GEN_16988 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10652 : rob_valid_28; // @[rob.scala 133:89 81:28]
  wire  _GEN_16989 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10653 : rob_valid_29; // @[rob.scala 133:89 81:28]
  wire  _GEN_16990 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10654 : rob_valid_30; // @[rob.scala 133:89 81:28]
  wire  _GEN_16991 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10655 : rob_valid_31; // @[rob.scala 133:89 81:28]
  wire  _GEN_16992 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10656 : rob_valid_32; // @[rob.scala 133:89 81:28]
  wire  _GEN_16993 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10657 : rob_valid_33; // @[rob.scala 133:89 81:28]
  wire  _GEN_16994 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10658 : rob_valid_34; // @[rob.scala 133:89 81:28]
  wire  _GEN_16995 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10659 : rob_valid_35; // @[rob.scala 133:89 81:28]
  wire  _GEN_16996 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10660 : rob_valid_36; // @[rob.scala 133:89 81:28]
  wire  _GEN_16997 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10661 : rob_valid_37; // @[rob.scala 133:89 81:28]
  wire  _GEN_16998 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10662 : rob_valid_38; // @[rob.scala 133:89 81:28]
  wire  _GEN_16999 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10663 : rob_valid_39; // @[rob.scala 133:89 81:28]
  wire  _GEN_17000 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10664 : rob_valid_40; // @[rob.scala 133:89 81:28]
  wire  _GEN_17001 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10665 : rob_valid_41; // @[rob.scala 133:89 81:28]
  wire  _GEN_17002 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10666 : rob_valid_42; // @[rob.scala 133:89 81:28]
  wire  _GEN_17003 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10667 : rob_valid_43; // @[rob.scala 133:89 81:28]
  wire  _GEN_17004 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10668 : rob_valid_44; // @[rob.scala 133:89 81:28]
  wire  _GEN_17005 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10669 : rob_valid_45; // @[rob.scala 133:89 81:28]
  wire  _GEN_17006 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10670 : rob_valid_46; // @[rob.scala 133:89 81:28]
  wire  _GEN_17007 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10671 : rob_valid_47; // @[rob.scala 133:89 81:28]
  wire  _GEN_17008 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10672 : rob_valid_48; // @[rob.scala 133:89 81:28]
  wire  _GEN_17009 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10673 : rob_valid_49; // @[rob.scala 133:89 81:28]
  wire  _GEN_17010 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10674 : rob_valid_50; // @[rob.scala 133:89 81:28]
  wire  _GEN_17011 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10675 : rob_valid_51; // @[rob.scala 133:89 81:28]
  wire  _GEN_17012 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10676 : rob_valid_52; // @[rob.scala 133:89 81:28]
  wire  _GEN_17013 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10677 : rob_valid_53; // @[rob.scala 133:89 81:28]
  wire  _GEN_17014 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10678 : rob_valid_54; // @[rob.scala 133:89 81:28]
  wire  _GEN_17015 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10679 : rob_valid_55; // @[rob.scala 133:89 81:28]
  wire  _GEN_17016 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10680 : rob_valid_56; // @[rob.scala 133:89 81:28]
  wire  _GEN_17017 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10681 : rob_valid_57; // @[rob.scala 133:89 81:28]
  wire  _GEN_17018 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10682 : rob_valid_58; // @[rob.scala 133:89 81:28]
  wire  _GEN_17019 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10683 : rob_valid_59; // @[rob.scala 133:89 81:28]
  wire  _GEN_17020 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10684 : rob_valid_60; // @[rob.scala 133:89 81:28]
  wire  _GEN_17021 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10685 : rob_valid_61; // @[rob.scala 133:89 81:28]
  wire  _GEN_17022 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10686 : rob_valid_62; // @[rob.scala 133:89 81:28]
  wire  _GEN_17023 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10687 : rob_valid_63; // @[rob.scala 133:89 81:28]
  wire [6:0] _GEN_17024 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _is_full_T_4 :
    allocate_ptr; // @[rob.scala 133:89 137:22 47:31]
  wire  _GEN_17025 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10688 : rob_done_0; // @[rob.scala 133:89 84:27]
  wire  _GEN_17026 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10689 : rob_done_1; // @[rob.scala 133:89 84:27]
  wire  _GEN_17027 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10690 : rob_done_2; // @[rob.scala 133:89 84:27]
  wire  _GEN_17028 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10691 : rob_done_3; // @[rob.scala 133:89 84:27]
  wire  _GEN_17029 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10692 : rob_done_4; // @[rob.scala 133:89 84:27]
  wire  _GEN_17030 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10693 : rob_done_5; // @[rob.scala 133:89 84:27]
  wire  _GEN_17031 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10694 : rob_done_6; // @[rob.scala 133:89 84:27]
  wire  _GEN_17032 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10695 : rob_done_7; // @[rob.scala 133:89 84:27]
  wire  _GEN_17033 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10696 : rob_done_8; // @[rob.scala 133:89 84:27]
  wire  _GEN_17034 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10697 : rob_done_9; // @[rob.scala 133:89 84:27]
  wire  _GEN_17035 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10698 : rob_done_10; // @[rob.scala 133:89 84:27]
  wire  _GEN_17036 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10699 : rob_done_11; // @[rob.scala 133:89 84:27]
  wire  _GEN_17037 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10700 : rob_done_12; // @[rob.scala 133:89 84:27]
  wire  _GEN_17038 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10701 : rob_done_13; // @[rob.scala 133:89 84:27]
  wire  _GEN_17039 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10702 : rob_done_14; // @[rob.scala 133:89 84:27]
  wire  _GEN_17040 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10703 : rob_done_15; // @[rob.scala 133:89 84:27]
  wire  _GEN_17041 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10704 : rob_done_16; // @[rob.scala 133:89 84:27]
  wire  _GEN_17042 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10705 : rob_done_17; // @[rob.scala 133:89 84:27]
  wire  _GEN_17043 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10706 : rob_done_18; // @[rob.scala 133:89 84:27]
  wire  _GEN_17044 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10707 : rob_done_19; // @[rob.scala 133:89 84:27]
  wire  _GEN_17045 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10708 : rob_done_20; // @[rob.scala 133:89 84:27]
  wire  _GEN_17046 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10709 : rob_done_21; // @[rob.scala 133:89 84:27]
  wire  _GEN_17047 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10710 : rob_done_22; // @[rob.scala 133:89 84:27]
  wire  _GEN_17048 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10711 : rob_done_23; // @[rob.scala 133:89 84:27]
  wire  _GEN_17049 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10712 : rob_done_24; // @[rob.scala 133:89 84:27]
  wire  _GEN_17050 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10713 : rob_done_25; // @[rob.scala 133:89 84:27]
  wire  _GEN_17051 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10714 : rob_done_26; // @[rob.scala 133:89 84:27]
  wire  _GEN_17052 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10715 : rob_done_27; // @[rob.scala 133:89 84:27]
  wire  _GEN_17053 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10716 : rob_done_28; // @[rob.scala 133:89 84:27]
  wire  _GEN_17054 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10717 : rob_done_29; // @[rob.scala 133:89 84:27]
  wire  _GEN_17055 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10718 : rob_done_30; // @[rob.scala 133:89 84:27]
  wire  _GEN_17056 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10719 : rob_done_31; // @[rob.scala 133:89 84:27]
  wire  _GEN_17057 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10720 : rob_done_32; // @[rob.scala 133:89 84:27]
  wire  _GEN_17058 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10721 : rob_done_33; // @[rob.scala 133:89 84:27]
  wire  _GEN_17059 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10722 : rob_done_34; // @[rob.scala 133:89 84:27]
  wire  _GEN_17060 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10723 : rob_done_35; // @[rob.scala 133:89 84:27]
  wire  _GEN_17061 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10724 : rob_done_36; // @[rob.scala 133:89 84:27]
  wire  _GEN_17062 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10725 : rob_done_37; // @[rob.scala 133:89 84:27]
  wire  _GEN_17063 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10726 : rob_done_38; // @[rob.scala 133:89 84:27]
  wire  _GEN_17064 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10727 : rob_done_39; // @[rob.scala 133:89 84:27]
  wire  _GEN_17065 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10728 : rob_done_40; // @[rob.scala 133:89 84:27]
  wire  _GEN_17066 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10729 : rob_done_41; // @[rob.scala 133:89 84:27]
  wire  _GEN_17067 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10730 : rob_done_42; // @[rob.scala 133:89 84:27]
  wire  _GEN_17068 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10731 : rob_done_43; // @[rob.scala 133:89 84:27]
  wire  _GEN_17069 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10732 : rob_done_44; // @[rob.scala 133:89 84:27]
  wire  _GEN_17070 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10733 : rob_done_45; // @[rob.scala 133:89 84:27]
  wire  _GEN_17071 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10734 : rob_done_46; // @[rob.scala 133:89 84:27]
  wire  _GEN_17072 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10735 : rob_done_47; // @[rob.scala 133:89 84:27]
  wire  _GEN_17073 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10736 : rob_done_48; // @[rob.scala 133:89 84:27]
  wire  _GEN_17074 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10737 : rob_done_49; // @[rob.scala 133:89 84:27]
  wire  _GEN_17075 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10738 : rob_done_50; // @[rob.scala 133:89 84:27]
  wire  _GEN_17076 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10739 : rob_done_51; // @[rob.scala 133:89 84:27]
  wire  _GEN_17077 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10740 : rob_done_52; // @[rob.scala 133:89 84:27]
  wire  _GEN_17078 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10741 : rob_done_53; // @[rob.scala 133:89 84:27]
  wire  _GEN_17079 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10742 : rob_done_54; // @[rob.scala 133:89 84:27]
  wire  _GEN_17080 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10743 : rob_done_55; // @[rob.scala 133:89 84:27]
  wire  _GEN_17081 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10744 : rob_done_56; // @[rob.scala 133:89 84:27]
  wire  _GEN_17082 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10745 : rob_done_57; // @[rob.scala 133:89 84:27]
  wire  _GEN_17083 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10746 : rob_done_58; // @[rob.scala 133:89 84:27]
  wire  _GEN_17084 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10747 : rob_done_59; // @[rob.scala 133:89 84:27]
  wire  _GEN_17085 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10748 : rob_done_60; // @[rob.scala 133:89 84:27]
  wire  _GEN_17086 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10749 : rob_done_61; // @[rob.scala 133:89 84:27]
  wire  _GEN_17087 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10750 : rob_done_62; // @[rob.scala 133:89 84:27]
  wire  _GEN_17088 = io_i_rob_allocation_reqs_0_valid | io_i_rob_allocation_reqs_1_valid ? _GEN_10751 : rob_done_63; // @[rob.scala 133:89 84:27]
  wire [31:0] _GEN_17153 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10816 : _GEN_15040
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17154 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10817 : _GEN_15041
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17155 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10818 : _GEN_15042
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17156 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10819 : _GEN_15043
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17157 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10820 : _GEN_15044
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17158 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10821 : _GEN_15045
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17159 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10822 : _GEN_15046
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17160 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10823 : _GEN_15047
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17161 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10824 : _GEN_15048
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17162 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10825 : _GEN_15049
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17163 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10826 : _GEN_15050
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17164 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10827 : _GEN_15051
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17165 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10828 : _GEN_15052
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17166 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10829 : _GEN_15053
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17167 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10830 : _GEN_15054
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17168 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10831 : _GEN_15055
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17169 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10832 : _GEN_15056
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17170 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10833 : _GEN_15057
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17171 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10834 : _GEN_15058
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17172 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10835 : _GEN_15059
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17173 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10836 : _GEN_15060
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17174 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10837 : _GEN_15061
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17175 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10838 : _GEN_15062
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17176 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10839 : _GEN_15063
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17177 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10840 : _GEN_15064
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17178 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10841 : _GEN_15065
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17179 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10842 : _GEN_15066
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17180 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10843 : _GEN_15067
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17181 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10844 : _GEN_15068
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17182 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10845 : _GEN_15069
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17183 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10846 : _GEN_15070
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17184 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10847 : _GEN_15071
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17185 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10848 : _GEN_15072
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17186 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10849 : _GEN_15073
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17187 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10850 : _GEN_15074
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17188 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10851 : _GEN_15075
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17189 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10852 : _GEN_15076
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17190 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10853 : _GEN_15077
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17191 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10854 : _GEN_15078
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17192 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10855 : _GEN_15079
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17193 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10856 : _GEN_15080
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17194 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10857 : _GEN_15081
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17195 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10858 : _GEN_15082
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17196 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10859 : _GEN_15083
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17197 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10860 : _GEN_15084
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17198 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10861 : _GEN_15085
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17199 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10862 : _GEN_15086
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17200 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10863 : _GEN_15087
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17201 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10864 : _GEN_15088
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17202 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10865 : _GEN_15089
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17203 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10866 : _GEN_15090
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17204 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10867 : _GEN_15091
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17205 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10868 : _GEN_15092
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17206 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10869 : _GEN_15093
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17207 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10870 : _GEN_15094
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17208 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10871 : _GEN_15095
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17209 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10872 : _GEN_15096
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17210 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10873 : _GEN_15097
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17211 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10874 : _GEN_15098
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17212 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10875 : _GEN_15099
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17213 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10876 : _GEN_15100
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17214 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10877 : _GEN_15101
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17215 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10878 : _GEN_15102
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17216 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10879 : _GEN_15103
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17217 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10880 : _GEN_15104
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17218 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10881 : _GEN_15105
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17219 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10882 : _GEN_15106
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17220 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10883 : _GEN_15107
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17221 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10884 : _GEN_15108
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17222 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10885 : _GEN_15109
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17223 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10886 : _GEN_15110
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17224 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10887 : _GEN_15111
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17225 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10888 : _GEN_15112
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17226 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10889 : _GEN_15113
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17227 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10890 : _GEN_15114
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17228 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10891 : _GEN_15115
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17229 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10892 : _GEN_15116
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17230 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10893 : _GEN_15117
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17231 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10894 : _GEN_15118
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17232 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10895 : _GEN_15119
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17233 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10896 : _GEN_15120
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17234 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10897 : _GEN_15121
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17235 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10898 : _GEN_15122
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17236 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10899 : _GEN_15123
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17237 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10900 : _GEN_15124
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17238 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10901 : _GEN_15125
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17239 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10902 : _GEN_15126
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17240 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10903 : _GEN_15127
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17241 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10904 : _GEN_15128
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17242 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10905 : _GEN_15129
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17243 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10906 : _GEN_15130
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17244 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10907 : _GEN_15131
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17245 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10908 : _GEN_15132
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17246 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10909 : _GEN_15133
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17247 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10910 : _GEN_15134
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17248 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10911 : _GEN_15135
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17249 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10912 : _GEN_15136
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17250 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10913 : _GEN_15137
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17251 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10914 : _GEN_15138
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17252 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10915 : _GEN_15139
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17253 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10916 : _GEN_15140
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17254 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10917 : _GEN_15141
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17255 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10918 : _GEN_15142
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17256 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10919 : _GEN_15143
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17257 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10920 : _GEN_15144
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17258 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10921 : _GEN_15145
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17259 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10922 : _GEN_15146
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17260 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10923 : _GEN_15147
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17261 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10924 : _GEN_15148
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17262 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10925 : _GEN_15149
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17263 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10926 : _GEN_15150
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17264 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10927 : _GEN_15151
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17265 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10928 : _GEN_15152
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17266 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10929 : _GEN_15153
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17267 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10930 : _GEN_15154
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17268 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10931 : _GEN_15155
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17269 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10932 : _GEN_15156
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17270 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10933 : _GEN_15157
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17271 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10934 : _GEN_15158
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17272 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10935 : _GEN_15159
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17273 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10936 : _GEN_15160
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17274 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10937 : _GEN_15161
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17275 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10938 : _GEN_15162
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17276 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10939 : _GEN_15163
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17277 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10940 : _GEN_15164
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17278 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10941 : _GEN_15165
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17279 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10942 : _GEN_15166
    ; // @[rob.scala 124:83]
  wire [31:0] _GEN_17280 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10943 : _GEN_15167
    ; // @[rob.scala 124:83]
  wire [6:0] _GEN_17281 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10944 : _GEN_15168; // @[rob.scala 124:83]
  wire [6:0] _GEN_17282 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10945 : _GEN_15169; // @[rob.scala 124:83]
  wire [6:0] _GEN_17283 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10946 : _GEN_15170; // @[rob.scala 124:83]
  wire [6:0] _GEN_17284 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10947 : _GEN_15171; // @[rob.scala 124:83]
  wire [6:0] _GEN_17285 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10948 : _GEN_15172; // @[rob.scala 124:83]
  wire [6:0] _GEN_17286 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10949 : _GEN_15173; // @[rob.scala 124:83]
  wire [6:0] _GEN_17287 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10950 : _GEN_15174; // @[rob.scala 124:83]
  wire [6:0] _GEN_17288 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10951 : _GEN_15175; // @[rob.scala 124:83]
  wire [6:0] _GEN_17289 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10952 : _GEN_15176; // @[rob.scala 124:83]
  wire [6:0] _GEN_17290 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10953 : _GEN_15177; // @[rob.scala 124:83]
  wire [6:0] _GEN_17291 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10954 : _GEN_15178; // @[rob.scala 124:83]
  wire [6:0] _GEN_17292 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10955 : _GEN_15179; // @[rob.scala 124:83]
  wire [6:0] _GEN_17293 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10956 : _GEN_15180; // @[rob.scala 124:83]
  wire [6:0] _GEN_17294 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10957 : _GEN_15181; // @[rob.scala 124:83]
  wire [6:0] _GEN_17295 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10958 : _GEN_15182; // @[rob.scala 124:83]
  wire [6:0] _GEN_17296 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10959 : _GEN_15183; // @[rob.scala 124:83]
  wire [6:0] _GEN_17297 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10960 : _GEN_15184; // @[rob.scala 124:83]
  wire [6:0] _GEN_17298 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10961 : _GEN_15185; // @[rob.scala 124:83]
  wire [6:0] _GEN_17299 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10962 : _GEN_15186; // @[rob.scala 124:83]
  wire [6:0] _GEN_17300 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10963 : _GEN_15187; // @[rob.scala 124:83]
  wire [6:0] _GEN_17301 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10964 : _GEN_15188; // @[rob.scala 124:83]
  wire [6:0] _GEN_17302 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10965 : _GEN_15189; // @[rob.scala 124:83]
  wire [6:0] _GEN_17303 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10966 : _GEN_15190; // @[rob.scala 124:83]
  wire [6:0] _GEN_17304 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10967 : _GEN_15191; // @[rob.scala 124:83]
  wire [6:0] _GEN_17305 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10968 : _GEN_15192; // @[rob.scala 124:83]
  wire [6:0] _GEN_17306 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10969 : _GEN_15193; // @[rob.scala 124:83]
  wire [6:0] _GEN_17307 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10970 : _GEN_15194; // @[rob.scala 124:83]
  wire [6:0] _GEN_17308 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10971 : _GEN_15195; // @[rob.scala 124:83]
  wire [6:0] _GEN_17309 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10972 : _GEN_15196; // @[rob.scala 124:83]
  wire [6:0] _GEN_17310 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10973 : _GEN_15197; // @[rob.scala 124:83]
  wire [6:0] _GEN_17311 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10974 : _GEN_15198; // @[rob.scala 124:83]
  wire [6:0] _GEN_17312 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10975 : _GEN_15199; // @[rob.scala 124:83]
  wire [6:0] _GEN_17313 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10976 : _GEN_15200; // @[rob.scala 124:83]
  wire [6:0] _GEN_17314 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10977 : _GEN_15201; // @[rob.scala 124:83]
  wire [6:0] _GEN_17315 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10978 : _GEN_15202; // @[rob.scala 124:83]
  wire [6:0] _GEN_17316 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10979 : _GEN_15203; // @[rob.scala 124:83]
  wire [6:0] _GEN_17317 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10980 : _GEN_15204; // @[rob.scala 124:83]
  wire [6:0] _GEN_17318 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10981 : _GEN_15205; // @[rob.scala 124:83]
  wire [6:0] _GEN_17319 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10982 : _GEN_15206; // @[rob.scala 124:83]
  wire [6:0] _GEN_17320 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10983 : _GEN_15207; // @[rob.scala 124:83]
  wire [6:0] _GEN_17321 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10984 : _GEN_15208; // @[rob.scala 124:83]
  wire [6:0] _GEN_17322 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10985 : _GEN_15209; // @[rob.scala 124:83]
  wire [6:0] _GEN_17323 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10986 : _GEN_15210; // @[rob.scala 124:83]
  wire [6:0] _GEN_17324 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10987 : _GEN_15211; // @[rob.scala 124:83]
  wire [6:0] _GEN_17325 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10988 : _GEN_15212; // @[rob.scala 124:83]
  wire [6:0] _GEN_17326 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10989 : _GEN_15213; // @[rob.scala 124:83]
  wire [6:0] _GEN_17327 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10990 : _GEN_15214; // @[rob.scala 124:83]
  wire [6:0] _GEN_17328 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10991 : _GEN_15215; // @[rob.scala 124:83]
  wire [6:0] _GEN_17329 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10992 : _GEN_15216; // @[rob.scala 124:83]
  wire [6:0] _GEN_17330 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10993 : _GEN_15217; // @[rob.scala 124:83]
  wire [6:0] _GEN_17331 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10994 : _GEN_15218; // @[rob.scala 124:83]
  wire [6:0] _GEN_17332 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10995 : _GEN_15219; // @[rob.scala 124:83]
  wire [6:0] _GEN_17333 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10996 : _GEN_15220; // @[rob.scala 124:83]
  wire [6:0] _GEN_17334 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10997 : _GEN_15221; // @[rob.scala 124:83]
  wire [6:0] _GEN_17335 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10998 : _GEN_15222; // @[rob.scala 124:83]
  wire [6:0] _GEN_17336 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_10999 : _GEN_15223; // @[rob.scala 124:83]
  wire [6:0] _GEN_17337 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11000 : _GEN_15224; // @[rob.scala 124:83]
  wire [6:0] _GEN_17338 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11001 : _GEN_15225; // @[rob.scala 124:83]
  wire [6:0] _GEN_17339 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11002 : _GEN_15226; // @[rob.scala 124:83]
  wire [6:0] _GEN_17340 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11003 : _GEN_15227; // @[rob.scala 124:83]
  wire [6:0] _GEN_17341 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11004 : _GEN_15228; // @[rob.scala 124:83]
  wire [6:0] _GEN_17342 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11005 : _GEN_15229; // @[rob.scala 124:83]
  wire [6:0] _GEN_17343 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11006 : _GEN_15230; // @[rob.scala 124:83]
  wire [6:0] _GEN_17344 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11007 : _GEN_15231; // @[rob.scala 124:83]
  wire [6:0] _GEN_17665 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11328 : _GEN_15552; // @[rob.scala 124:83]
  wire [6:0] _GEN_17666 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11329 : _GEN_15553; // @[rob.scala 124:83]
  wire [6:0] _GEN_17667 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11330 : _GEN_15554; // @[rob.scala 124:83]
  wire [6:0] _GEN_17668 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11331 : _GEN_15555; // @[rob.scala 124:83]
  wire [6:0] _GEN_17669 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11332 : _GEN_15556; // @[rob.scala 124:83]
  wire [6:0] _GEN_17670 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11333 : _GEN_15557; // @[rob.scala 124:83]
  wire [6:0] _GEN_17671 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11334 : _GEN_15558; // @[rob.scala 124:83]
  wire [6:0] _GEN_17672 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11335 : _GEN_15559; // @[rob.scala 124:83]
  wire [6:0] _GEN_17673 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11336 : _GEN_15560; // @[rob.scala 124:83]
  wire [6:0] _GEN_17674 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11337 : _GEN_15561; // @[rob.scala 124:83]
  wire [6:0] _GEN_17675 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11338 : _GEN_15562; // @[rob.scala 124:83]
  wire [6:0] _GEN_17676 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11339 : _GEN_15563; // @[rob.scala 124:83]
  wire [6:0] _GEN_17677 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11340 : _GEN_15564; // @[rob.scala 124:83]
  wire [6:0] _GEN_17678 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11341 : _GEN_15565; // @[rob.scala 124:83]
  wire [6:0] _GEN_17679 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11342 : _GEN_15566; // @[rob.scala 124:83]
  wire [6:0] _GEN_17680 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11343 : _GEN_15567; // @[rob.scala 124:83]
  wire [6:0] _GEN_17681 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11344 : _GEN_15568; // @[rob.scala 124:83]
  wire [6:0] _GEN_17682 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11345 : _GEN_15569; // @[rob.scala 124:83]
  wire [6:0] _GEN_17683 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11346 : _GEN_15570; // @[rob.scala 124:83]
  wire [6:0] _GEN_17684 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11347 : _GEN_15571; // @[rob.scala 124:83]
  wire [6:0] _GEN_17685 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11348 : _GEN_15572; // @[rob.scala 124:83]
  wire [6:0] _GEN_17686 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11349 : _GEN_15573; // @[rob.scala 124:83]
  wire [6:0] _GEN_17687 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11350 : _GEN_15574; // @[rob.scala 124:83]
  wire [6:0] _GEN_17688 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11351 : _GEN_15575; // @[rob.scala 124:83]
  wire [6:0] _GEN_17689 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11352 : _GEN_15576; // @[rob.scala 124:83]
  wire [6:0] _GEN_17690 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11353 : _GEN_15577; // @[rob.scala 124:83]
  wire [6:0] _GEN_17691 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11354 : _GEN_15578; // @[rob.scala 124:83]
  wire [6:0] _GEN_17692 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11355 : _GEN_15579; // @[rob.scala 124:83]
  wire [6:0] _GEN_17693 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11356 : _GEN_15580; // @[rob.scala 124:83]
  wire [6:0] _GEN_17694 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11357 : _GEN_15581; // @[rob.scala 124:83]
  wire [6:0] _GEN_17695 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11358 : _GEN_15582; // @[rob.scala 124:83]
  wire [6:0] _GEN_17696 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11359 : _GEN_15583; // @[rob.scala 124:83]
  wire [6:0] _GEN_17697 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11360 : _GEN_15584; // @[rob.scala 124:83]
  wire [6:0] _GEN_17698 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11361 : _GEN_15585; // @[rob.scala 124:83]
  wire [6:0] _GEN_17699 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11362 : _GEN_15586; // @[rob.scala 124:83]
  wire [6:0] _GEN_17700 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11363 : _GEN_15587; // @[rob.scala 124:83]
  wire [6:0] _GEN_17701 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11364 : _GEN_15588; // @[rob.scala 124:83]
  wire [6:0] _GEN_17702 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11365 : _GEN_15589; // @[rob.scala 124:83]
  wire [6:0] _GEN_17703 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11366 : _GEN_15590; // @[rob.scala 124:83]
  wire [6:0] _GEN_17704 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11367 : _GEN_15591; // @[rob.scala 124:83]
  wire [6:0] _GEN_17705 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11368 : _GEN_15592; // @[rob.scala 124:83]
  wire [6:0] _GEN_17706 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11369 : _GEN_15593; // @[rob.scala 124:83]
  wire [6:0] _GEN_17707 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11370 : _GEN_15594; // @[rob.scala 124:83]
  wire [6:0] _GEN_17708 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11371 : _GEN_15595; // @[rob.scala 124:83]
  wire [6:0] _GEN_17709 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11372 : _GEN_15596; // @[rob.scala 124:83]
  wire [6:0] _GEN_17710 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11373 : _GEN_15597; // @[rob.scala 124:83]
  wire [6:0] _GEN_17711 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11374 : _GEN_15598; // @[rob.scala 124:83]
  wire [6:0] _GEN_17712 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11375 : _GEN_15599; // @[rob.scala 124:83]
  wire [6:0] _GEN_17713 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11376 : _GEN_15600; // @[rob.scala 124:83]
  wire [6:0] _GEN_17714 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11377 : _GEN_15601; // @[rob.scala 124:83]
  wire [6:0] _GEN_17715 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11378 : _GEN_15602; // @[rob.scala 124:83]
  wire [6:0] _GEN_17716 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11379 : _GEN_15603; // @[rob.scala 124:83]
  wire [6:0] _GEN_17717 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11380 : _GEN_15604; // @[rob.scala 124:83]
  wire [6:0] _GEN_17718 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11381 : _GEN_15605; // @[rob.scala 124:83]
  wire [6:0] _GEN_17719 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11382 : _GEN_15606; // @[rob.scala 124:83]
  wire [6:0] _GEN_17720 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11383 : _GEN_15607; // @[rob.scala 124:83]
  wire [6:0] _GEN_17721 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11384 : _GEN_15608; // @[rob.scala 124:83]
  wire [6:0] _GEN_17722 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11385 : _GEN_15609; // @[rob.scala 124:83]
  wire [6:0] _GEN_17723 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11386 : _GEN_15610; // @[rob.scala 124:83]
  wire [6:0] _GEN_17724 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11387 : _GEN_15611; // @[rob.scala 124:83]
  wire [6:0] _GEN_17725 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11388 : _GEN_15612; // @[rob.scala 124:83]
  wire [6:0] _GEN_17726 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11389 : _GEN_15613; // @[rob.scala 124:83]
  wire [6:0] _GEN_17727 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11390 : _GEN_15614; // @[rob.scala 124:83]
  wire [6:0] _GEN_17728 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11391 : _GEN_15615; // @[rob.scala 124:83]
  wire [6:0] _GEN_17729 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11392 : _GEN_15616; // @[rob.scala 124:83]
  wire [6:0] _GEN_17730 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11393 : _GEN_15617; // @[rob.scala 124:83]
  wire [6:0] _GEN_17731 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11394 : _GEN_15618; // @[rob.scala 124:83]
  wire [6:0] _GEN_17732 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11395 : _GEN_15619; // @[rob.scala 124:83]
  wire [6:0] _GEN_17733 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11396 : _GEN_15620; // @[rob.scala 124:83]
  wire [6:0] _GEN_17734 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11397 : _GEN_15621; // @[rob.scala 124:83]
  wire [6:0] _GEN_17735 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11398 : _GEN_15622; // @[rob.scala 124:83]
  wire [6:0] _GEN_17736 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11399 : _GEN_15623; // @[rob.scala 124:83]
  wire [6:0] _GEN_17737 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11400 : _GEN_15624; // @[rob.scala 124:83]
  wire [6:0] _GEN_17738 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11401 : _GEN_15625; // @[rob.scala 124:83]
  wire [6:0] _GEN_17739 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11402 : _GEN_15626; // @[rob.scala 124:83]
  wire [6:0] _GEN_17740 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11403 : _GEN_15627; // @[rob.scala 124:83]
  wire [6:0] _GEN_17741 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11404 : _GEN_15628; // @[rob.scala 124:83]
  wire [6:0] _GEN_17742 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11405 : _GEN_15629; // @[rob.scala 124:83]
  wire [6:0] _GEN_17743 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11406 : _GEN_15630; // @[rob.scala 124:83]
  wire [6:0] _GEN_17744 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11407 : _GEN_15631; // @[rob.scala 124:83]
  wire [6:0] _GEN_17745 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11408 : _GEN_15632; // @[rob.scala 124:83]
  wire [6:0] _GEN_17746 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11409 : _GEN_15633; // @[rob.scala 124:83]
  wire [6:0] _GEN_17747 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11410 : _GEN_15634; // @[rob.scala 124:83]
  wire [6:0] _GEN_17748 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11411 : _GEN_15635; // @[rob.scala 124:83]
  wire [6:0] _GEN_17749 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11412 : _GEN_15636; // @[rob.scala 124:83]
  wire [6:0] _GEN_17750 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11413 : _GEN_15637; // @[rob.scala 124:83]
  wire [6:0] _GEN_17751 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11414 : _GEN_15638; // @[rob.scala 124:83]
  wire [6:0] _GEN_17752 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11415 : _GEN_15639; // @[rob.scala 124:83]
  wire [6:0] _GEN_17753 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11416 : _GEN_15640; // @[rob.scala 124:83]
  wire [6:0] _GEN_17754 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11417 : _GEN_15641; // @[rob.scala 124:83]
  wire [6:0] _GEN_17755 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11418 : _GEN_15642; // @[rob.scala 124:83]
  wire [6:0] _GEN_17756 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11419 : _GEN_15643; // @[rob.scala 124:83]
  wire [6:0] _GEN_17757 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11420 : _GEN_15644; // @[rob.scala 124:83]
  wire [6:0] _GEN_17758 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11421 : _GEN_15645; // @[rob.scala 124:83]
  wire [6:0] _GEN_17759 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11422 : _GEN_15646; // @[rob.scala 124:83]
  wire [6:0] _GEN_17760 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11423 : _GEN_15647; // @[rob.scala 124:83]
  wire [6:0] _GEN_17761 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11424 : _GEN_15648; // @[rob.scala 124:83]
  wire [6:0] _GEN_17762 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11425 : _GEN_15649; // @[rob.scala 124:83]
  wire [6:0] _GEN_17763 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11426 : _GEN_15650; // @[rob.scala 124:83]
  wire [6:0] _GEN_17764 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11427 : _GEN_15651; // @[rob.scala 124:83]
  wire [6:0] _GEN_17765 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11428 : _GEN_15652; // @[rob.scala 124:83]
  wire [6:0] _GEN_17766 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11429 : _GEN_15653; // @[rob.scala 124:83]
  wire [6:0] _GEN_17767 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11430 : _GEN_15654; // @[rob.scala 124:83]
  wire [6:0] _GEN_17768 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11431 : _GEN_15655; // @[rob.scala 124:83]
  wire [6:0] _GEN_17769 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11432 : _GEN_15656; // @[rob.scala 124:83]
  wire [6:0] _GEN_17770 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11433 : _GEN_15657; // @[rob.scala 124:83]
  wire [6:0] _GEN_17771 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11434 : _GEN_15658; // @[rob.scala 124:83]
  wire [6:0] _GEN_17772 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11435 : _GEN_15659; // @[rob.scala 124:83]
  wire [6:0] _GEN_17773 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11436 : _GEN_15660; // @[rob.scala 124:83]
  wire [6:0] _GEN_17774 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11437 : _GEN_15661; // @[rob.scala 124:83]
  wire [6:0] _GEN_17775 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11438 : _GEN_15662; // @[rob.scala 124:83]
  wire [6:0] _GEN_17776 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11439 : _GEN_15663; // @[rob.scala 124:83]
  wire [6:0] _GEN_17777 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11440 : _GEN_15664; // @[rob.scala 124:83]
  wire [6:0] _GEN_17778 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11441 : _GEN_15665; // @[rob.scala 124:83]
  wire [6:0] _GEN_17779 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11442 : _GEN_15666; // @[rob.scala 124:83]
  wire [6:0] _GEN_17780 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11443 : _GEN_15667; // @[rob.scala 124:83]
  wire [6:0] _GEN_17781 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11444 : _GEN_15668; // @[rob.scala 124:83]
  wire [6:0] _GEN_17782 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11445 : _GEN_15669; // @[rob.scala 124:83]
  wire [6:0] _GEN_17783 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11446 : _GEN_15670; // @[rob.scala 124:83]
  wire [6:0] _GEN_17784 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11447 : _GEN_15671; // @[rob.scala 124:83]
  wire [6:0] _GEN_17785 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11448 : _GEN_15672; // @[rob.scala 124:83]
  wire [6:0] _GEN_17786 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11449 : _GEN_15673; // @[rob.scala 124:83]
  wire [6:0] _GEN_17787 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11450 : _GEN_15674; // @[rob.scala 124:83]
  wire [6:0] _GEN_17788 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11451 : _GEN_15675; // @[rob.scala 124:83]
  wire [6:0] _GEN_17789 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11452 : _GEN_15676; // @[rob.scala 124:83]
  wire [6:0] _GEN_17790 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11453 : _GEN_15677; // @[rob.scala 124:83]
  wire [6:0] _GEN_17791 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11454 : _GEN_15678; // @[rob.scala 124:83]
  wire [6:0] _GEN_17792 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11455 : _GEN_15679; // @[rob.scala 124:83]
  wire [4:0] _GEN_17793 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11456 : _GEN_15680; // @[rob.scala 124:83]
  wire [4:0] _GEN_17794 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11457 : _GEN_15681; // @[rob.scala 124:83]
  wire [4:0] _GEN_17795 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11458 : _GEN_15682; // @[rob.scala 124:83]
  wire [4:0] _GEN_17796 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11459 : _GEN_15683; // @[rob.scala 124:83]
  wire [4:0] _GEN_17797 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11460 : _GEN_15684; // @[rob.scala 124:83]
  wire [4:0] _GEN_17798 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11461 : _GEN_15685; // @[rob.scala 124:83]
  wire [4:0] _GEN_17799 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11462 : _GEN_15686; // @[rob.scala 124:83]
  wire [4:0] _GEN_17800 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11463 : _GEN_15687; // @[rob.scala 124:83]
  wire [4:0] _GEN_17801 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11464 : _GEN_15688; // @[rob.scala 124:83]
  wire [4:0] _GEN_17802 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11465 : _GEN_15689; // @[rob.scala 124:83]
  wire [4:0] _GEN_17803 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11466 : _GEN_15690; // @[rob.scala 124:83]
  wire [4:0] _GEN_17804 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11467 : _GEN_15691; // @[rob.scala 124:83]
  wire [4:0] _GEN_17805 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11468 : _GEN_15692; // @[rob.scala 124:83]
  wire [4:0] _GEN_17806 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11469 : _GEN_15693; // @[rob.scala 124:83]
  wire [4:0] _GEN_17807 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11470 : _GEN_15694; // @[rob.scala 124:83]
  wire [4:0] _GEN_17808 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11471 : _GEN_15695; // @[rob.scala 124:83]
  wire [4:0] _GEN_17809 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11472 : _GEN_15696; // @[rob.scala 124:83]
  wire [4:0] _GEN_17810 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11473 : _GEN_15697; // @[rob.scala 124:83]
  wire [4:0] _GEN_17811 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11474 : _GEN_15698; // @[rob.scala 124:83]
  wire [4:0] _GEN_17812 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11475 : _GEN_15699; // @[rob.scala 124:83]
  wire [4:0] _GEN_17813 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11476 : _GEN_15700; // @[rob.scala 124:83]
  wire [4:0] _GEN_17814 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11477 : _GEN_15701; // @[rob.scala 124:83]
  wire [4:0] _GEN_17815 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11478 : _GEN_15702; // @[rob.scala 124:83]
  wire [4:0] _GEN_17816 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11479 : _GEN_15703; // @[rob.scala 124:83]
  wire [4:0] _GEN_17817 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11480 : _GEN_15704; // @[rob.scala 124:83]
  wire [4:0] _GEN_17818 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11481 : _GEN_15705; // @[rob.scala 124:83]
  wire [4:0] _GEN_17819 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11482 : _GEN_15706; // @[rob.scala 124:83]
  wire [4:0] _GEN_17820 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11483 : _GEN_15707; // @[rob.scala 124:83]
  wire [4:0] _GEN_17821 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11484 : _GEN_15708; // @[rob.scala 124:83]
  wire [4:0] _GEN_17822 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11485 : _GEN_15709; // @[rob.scala 124:83]
  wire [4:0] _GEN_17823 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11486 : _GEN_15710; // @[rob.scala 124:83]
  wire [4:0] _GEN_17824 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11487 : _GEN_15711; // @[rob.scala 124:83]
  wire [4:0] _GEN_17825 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11488 : _GEN_15712; // @[rob.scala 124:83]
  wire [4:0] _GEN_17826 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11489 : _GEN_15713; // @[rob.scala 124:83]
  wire [4:0] _GEN_17827 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11490 : _GEN_15714; // @[rob.scala 124:83]
  wire [4:0] _GEN_17828 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11491 : _GEN_15715; // @[rob.scala 124:83]
  wire [4:0] _GEN_17829 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11492 : _GEN_15716; // @[rob.scala 124:83]
  wire [4:0] _GEN_17830 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11493 : _GEN_15717; // @[rob.scala 124:83]
  wire [4:0] _GEN_17831 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11494 : _GEN_15718; // @[rob.scala 124:83]
  wire [4:0] _GEN_17832 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11495 : _GEN_15719; // @[rob.scala 124:83]
  wire [4:0] _GEN_17833 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11496 : _GEN_15720; // @[rob.scala 124:83]
  wire [4:0] _GEN_17834 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11497 : _GEN_15721; // @[rob.scala 124:83]
  wire [4:0] _GEN_17835 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11498 : _GEN_15722; // @[rob.scala 124:83]
  wire [4:0] _GEN_17836 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11499 : _GEN_15723; // @[rob.scala 124:83]
  wire [4:0] _GEN_17837 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11500 : _GEN_15724; // @[rob.scala 124:83]
  wire [4:0] _GEN_17838 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11501 : _GEN_15725; // @[rob.scala 124:83]
  wire [4:0] _GEN_17839 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11502 : _GEN_15726; // @[rob.scala 124:83]
  wire [4:0] _GEN_17840 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11503 : _GEN_15727; // @[rob.scala 124:83]
  wire [4:0] _GEN_17841 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11504 : _GEN_15728; // @[rob.scala 124:83]
  wire [4:0] _GEN_17842 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11505 : _GEN_15729; // @[rob.scala 124:83]
  wire [4:0] _GEN_17843 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11506 : _GEN_15730; // @[rob.scala 124:83]
  wire [4:0] _GEN_17844 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11507 : _GEN_15731; // @[rob.scala 124:83]
  wire [4:0] _GEN_17845 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11508 : _GEN_15732; // @[rob.scala 124:83]
  wire [4:0] _GEN_17846 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11509 : _GEN_15733; // @[rob.scala 124:83]
  wire [4:0] _GEN_17847 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11510 : _GEN_15734; // @[rob.scala 124:83]
  wire [4:0] _GEN_17848 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11511 : _GEN_15735; // @[rob.scala 124:83]
  wire [4:0] _GEN_17849 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11512 : _GEN_15736; // @[rob.scala 124:83]
  wire [4:0] _GEN_17850 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11513 : _GEN_15737; // @[rob.scala 124:83]
  wire [4:0] _GEN_17851 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11514 : _GEN_15738; // @[rob.scala 124:83]
  wire [4:0] _GEN_17852 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11515 : _GEN_15739; // @[rob.scala 124:83]
  wire [4:0] _GEN_17853 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11516 : _GEN_15740; // @[rob.scala 124:83]
  wire [4:0] _GEN_17854 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11517 : _GEN_15741; // @[rob.scala 124:83]
  wire [4:0] _GEN_17855 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11518 : _GEN_15742; // @[rob.scala 124:83]
  wire [4:0] _GEN_17856 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_11519 : _GEN_15743; // @[rob.scala 124:83]
  wire [63:0] _GEN_18497 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12160 : _GEN_16384
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18498 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12161 : _GEN_16385
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18499 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12162 : _GEN_16386
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18500 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12163 : _GEN_16387
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18501 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12164 : _GEN_16388
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18502 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12165 : _GEN_16389
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18503 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12166 : _GEN_16390
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18504 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12167 : _GEN_16391
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18505 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12168 : _GEN_16392
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18506 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12169 : _GEN_16393
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18507 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12170 : _GEN_16394
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18508 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12171 : _GEN_16395
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18509 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12172 : _GEN_16396
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18510 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12173 : _GEN_16397
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18511 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12174 : _GEN_16398
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18512 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12175 : _GEN_16399
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18513 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12176 : _GEN_16400
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18514 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12177 : _GEN_16401
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18515 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12178 : _GEN_16402
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18516 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12179 : _GEN_16403
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18517 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12180 : _GEN_16404
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18518 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12181 : _GEN_16405
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18519 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12182 : _GEN_16406
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18520 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12183 : _GEN_16407
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18521 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12184 : _GEN_16408
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18522 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12185 : _GEN_16409
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18523 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12186 : _GEN_16410
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18524 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12187 : _GEN_16411
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18525 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12188 : _GEN_16412
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18526 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12189 : _GEN_16413
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18527 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12190 : _GEN_16414
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18528 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12191 : _GEN_16415
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18529 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12192 : _GEN_16416
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18530 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12193 : _GEN_16417
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18531 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12194 : _GEN_16418
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18532 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12195 : _GEN_16419
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18533 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12196 : _GEN_16420
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18534 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12197 : _GEN_16421
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18535 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12198 : _GEN_16422
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18536 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12199 : _GEN_16423
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18537 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12200 : _GEN_16424
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18538 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12201 : _GEN_16425
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18539 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12202 : _GEN_16426
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18540 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12203 : _GEN_16427
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18541 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12204 : _GEN_16428
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18542 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12205 : _GEN_16429
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18543 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12206 : _GEN_16430
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18544 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12207 : _GEN_16431
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18545 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12208 : _GEN_16432
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18546 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12209 : _GEN_16433
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18547 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12210 : _GEN_16434
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18548 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12211 : _GEN_16435
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18549 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12212 : _GEN_16436
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18550 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12213 : _GEN_16437
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18551 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12214 : _GEN_16438
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18552 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12215 : _GEN_16439
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18553 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12216 : _GEN_16440
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18554 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12217 : _GEN_16441
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18555 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12218 : _GEN_16442
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18556 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12219 : _GEN_16443
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18557 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12220 : _GEN_16444
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18558 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12221 : _GEN_16445
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18559 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12222 : _GEN_16446
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18560 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12223 : _GEN_16447
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18561 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12224 : _GEN_16448
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18562 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12225 : _GEN_16449
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18563 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12226 : _GEN_16450
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18564 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12227 : _GEN_16451
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18565 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12228 : _GEN_16452
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18566 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12229 : _GEN_16453
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18567 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12230 : _GEN_16454
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18568 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12231 : _GEN_16455
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18569 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12232 : _GEN_16456
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18570 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12233 : _GEN_16457
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18571 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12234 : _GEN_16458
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18572 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12235 : _GEN_16459
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18573 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12236 : _GEN_16460
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18574 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12237 : _GEN_16461
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18575 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12238 : _GEN_16462
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18576 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12239 : _GEN_16463
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18577 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12240 : _GEN_16464
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18578 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12241 : _GEN_16465
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18579 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12242 : _GEN_16466
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18580 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12243 : _GEN_16467
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18581 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12244 : _GEN_16468
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18582 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12245 : _GEN_16469
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18583 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12246 : _GEN_16470
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18584 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12247 : _GEN_16471
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18585 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12248 : _GEN_16472
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18586 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12249 : _GEN_16473
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18587 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12250 : _GEN_16474
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18588 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12251 : _GEN_16475
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18589 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12252 : _GEN_16476
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18590 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12253 : _GEN_16477
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18591 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12254 : _GEN_16478
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18592 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12255 : _GEN_16479
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18593 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12256 : _GEN_16480
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18594 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12257 : _GEN_16481
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18595 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12258 : _GEN_16482
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18596 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12259 : _GEN_16483
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18597 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12260 : _GEN_16484
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18598 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12261 : _GEN_16485
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18599 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12262 : _GEN_16486
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18600 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12263 : _GEN_16487
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18601 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12264 : _GEN_16488
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18602 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12265 : _GEN_16489
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18603 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12266 : _GEN_16490
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18604 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12267 : _GEN_16491
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18605 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12268 : _GEN_16492
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18606 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12269 : _GEN_16493
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18607 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12270 : _GEN_16494
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18608 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12271 : _GEN_16495
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18609 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12272 : _GEN_16496
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18610 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12273 : _GEN_16497
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18611 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12274 : _GEN_16498
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18612 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12275 : _GEN_16499
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18613 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12276 : _GEN_16500
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18614 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12277 : _GEN_16501
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18615 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12278 : _GEN_16502
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18616 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12279 : _GEN_16503
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18617 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12280 : _GEN_16504
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18618 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12281 : _GEN_16505
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18619 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12282 : _GEN_16506
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18620 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12283 : _GEN_16507
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18621 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12284 : _GEN_16508
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18622 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12285 : _GEN_16509
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18623 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12286 : _GEN_16510
    ; // @[rob.scala 124:83]
  wire [63:0] _GEN_18624 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12287 : _GEN_16511
    ; // @[rob.scala 124:83]
  wire [4:0] _GEN_18881 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12544 : _GEN_16768; // @[rob.scala 124:83]
  wire [4:0] _GEN_18882 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12545 : _GEN_16769; // @[rob.scala 124:83]
  wire [4:0] _GEN_18883 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12546 : _GEN_16770; // @[rob.scala 124:83]
  wire [4:0] _GEN_18884 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12547 : _GEN_16771; // @[rob.scala 124:83]
  wire [4:0] _GEN_18885 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12548 : _GEN_16772; // @[rob.scala 124:83]
  wire [4:0] _GEN_18886 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12549 : _GEN_16773; // @[rob.scala 124:83]
  wire [4:0] _GEN_18887 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12550 : _GEN_16774; // @[rob.scala 124:83]
  wire [4:0] _GEN_18888 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12551 : _GEN_16775; // @[rob.scala 124:83]
  wire [4:0] _GEN_18889 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12552 : _GEN_16776; // @[rob.scala 124:83]
  wire [4:0] _GEN_18890 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12553 : _GEN_16777; // @[rob.scala 124:83]
  wire [4:0] _GEN_18891 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12554 : _GEN_16778; // @[rob.scala 124:83]
  wire [4:0] _GEN_18892 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12555 : _GEN_16779; // @[rob.scala 124:83]
  wire [4:0] _GEN_18893 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12556 : _GEN_16780; // @[rob.scala 124:83]
  wire [4:0] _GEN_18894 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12557 : _GEN_16781; // @[rob.scala 124:83]
  wire [4:0] _GEN_18895 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12558 : _GEN_16782; // @[rob.scala 124:83]
  wire [4:0] _GEN_18896 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12559 : _GEN_16783; // @[rob.scala 124:83]
  wire [4:0] _GEN_18897 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12560 : _GEN_16784; // @[rob.scala 124:83]
  wire [4:0] _GEN_18898 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12561 : _GEN_16785; // @[rob.scala 124:83]
  wire [4:0] _GEN_18899 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12562 : _GEN_16786; // @[rob.scala 124:83]
  wire [4:0] _GEN_18900 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12563 : _GEN_16787; // @[rob.scala 124:83]
  wire [4:0] _GEN_18901 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12564 : _GEN_16788; // @[rob.scala 124:83]
  wire [4:0] _GEN_18902 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12565 : _GEN_16789; // @[rob.scala 124:83]
  wire [4:0] _GEN_18903 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12566 : _GEN_16790; // @[rob.scala 124:83]
  wire [4:0] _GEN_18904 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12567 : _GEN_16791; // @[rob.scala 124:83]
  wire [4:0] _GEN_18905 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12568 : _GEN_16792; // @[rob.scala 124:83]
  wire [4:0] _GEN_18906 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12569 : _GEN_16793; // @[rob.scala 124:83]
  wire [4:0] _GEN_18907 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12570 : _GEN_16794; // @[rob.scala 124:83]
  wire [4:0] _GEN_18908 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12571 : _GEN_16795; // @[rob.scala 124:83]
  wire [4:0] _GEN_18909 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12572 : _GEN_16796; // @[rob.scala 124:83]
  wire [4:0] _GEN_18910 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12573 : _GEN_16797; // @[rob.scala 124:83]
  wire [4:0] _GEN_18911 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12574 : _GEN_16798; // @[rob.scala 124:83]
  wire [4:0] _GEN_18912 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12575 : _GEN_16799; // @[rob.scala 124:83]
  wire [4:0] _GEN_18913 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12576 : _GEN_16800; // @[rob.scala 124:83]
  wire [4:0] _GEN_18914 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12577 : _GEN_16801; // @[rob.scala 124:83]
  wire [4:0] _GEN_18915 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12578 : _GEN_16802; // @[rob.scala 124:83]
  wire [4:0] _GEN_18916 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12579 : _GEN_16803; // @[rob.scala 124:83]
  wire [4:0] _GEN_18917 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12580 : _GEN_16804; // @[rob.scala 124:83]
  wire [4:0] _GEN_18918 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12581 : _GEN_16805; // @[rob.scala 124:83]
  wire [4:0] _GEN_18919 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12582 : _GEN_16806; // @[rob.scala 124:83]
  wire [4:0] _GEN_18920 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12583 : _GEN_16807; // @[rob.scala 124:83]
  wire [4:0] _GEN_18921 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12584 : _GEN_16808; // @[rob.scala 124:83]
  wire [4:0] _GEN_18922 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12585 : _GEN_16809; // @[rob.scala 124:83]
  wire [4:0] _GEN_18923 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12586 : _GEN_16810; // @[rob.scala 124:83]
  wire [4:0] _GEN_18924 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12587 : _GEN_16811; // @[rob.scala 124:83]
  wire [4:0] _GEN_18925 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12588 : _GEN_16812; // @[rob.scala 124:83]
  wire [4:0] _GEN_18926 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12589 : _GEN_16813; // @[rob.scala 124:83]
  wire [4:0] _GEN_18927 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12590 : _GEN_16814; // @[rob.scala 124:83]
  wire [4:0] _GEN_18928 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12591 : _GEN_16815; // @[rob.scala 124:83]
  wire [4:0] _GEN_18929 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12592 : _GEN_16816; // @[rob.scala 124:83]
  wire [4:0] _GEN_18930 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12593 : _GEN_16817; // @[rob.scala 124:83]
  wire [4:0] _GEN_18931 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12594 : _GEN_16818; // @[rob.scala 124:83]
  wire [4:0] _GEN_18932 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12595 : _GEN_16819; // @[rob.scala 124:83]
  wire [4:0] _GEN_18933 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12596 : _GEN_16820; // @[rob.scala 124:83]
  wire [4:0] _GEN_18934 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12597 : _GEN_16821; // @[rob.scala 124:83]
  wire [4:0] _GEN_18935 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12598 : _GEN_16822; // @[rob.scala 124:83]
  wire [4:0] _GEN_18936 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12599 : _GEN_16823; // @[rob.scala 124:83]
  wire [4:0] _GEN_18937 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12600 : _GEN_16824; // @[rob.scala 124:83]
  wire [4:0] _GEN_18938 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12601 : _GEN_16825; // @[rob.scala 124:83]
  wire [4:0] _GEN_18939 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12602 : _GEN_16826; // @[rob.scala 124:83]
  wire [4:0] _GEN_18940 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12603 : _GEN_16827; // @[rob.scala 124:83]
  wire [4:0] _GEN_18941 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12604 : _GEN_16828; // @[rob.scala 124:83]
  wire [4:0] _GEN_18942 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12605 : _GEN_16829; // @[rob.scala 124:83]
  wire [4:0] _GEN_18943 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12606 : _GEN_16830; // @[rob.scala 124:83]
  wire [4:0] _GEN_18944 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12607 : _GEN_16831; // @[rob.scala 124:83]
  wire  _GEN_19073 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12736 : _GEN_16960; // @[rob.scala 124:83]
  wire  _GEN_19074 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12737 : _GEN_16961; // @[rob.scala 124:83]
  wire  _GEN_19075 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12738 : _GEN_16962; // @[rob.scala 124:83]
  wire  _GEN_19076 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12739 : _GEN_16963; // @[rob.scala 124:83]
  wire  _GEN_19077 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12740 : _GEN_16964; // @[rob.scala 124:83]
  wire  _GEN_19078 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12741 : _GEN_16965; // @[rob.scala 124:83]
  wire  _GEN_19079 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12742 : _GEN_16966; // @[rob.scala 124:83]
  wire  _GEN_19080 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12743 : _GEN_16967; // @[rob.scala 124:83]
  wire  _GEN_19081 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12744 : _GEN_16968; // @[rob.scala 124:83]
  wire  _GEN_19082 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12745 : _GEN_16969; // @[rob.scala 124:83]
  wire  _GEN_19083 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12746 : _GEN_16970; // @[rob.scala 124:83]
  wire  _GEN_19084 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12747 : _GEN_16971; // @[rob.scala 124:83]
  wire  _GEN_19085 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12748 : _GEN_16972; // @[rob.scala 124:83]
  wire  _GEN_19086 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12749 : _GEN_16973; // @[rob.scala 124:83]
  wire  _GEN_19087 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12750 : _GEN_16974; // @[rob.scala 124:83]
  wire  _GEN_19088 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12751 : _GEN_16975; // @[rob.scala 124:83]
  wire  _GEN_19089 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12752 : _GEN_16976; // @[rob.scala 124:83]
  wire  _GEN_19090 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12753 : _GEN_16977; // @[rob.scala 124:83]
  wire  _GEN_19091 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12754 : _GEN_16978; // @[rob.scala 124:83]
  wire  _GEN_19092 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12755 : _GEN_16979; // @[rob.scala 124:83]
  wire  _GEN_19093 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12756 : _GEN_16980; // @[rob.scala 124:83]
  wire  _GEN_19094 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12757 : _GEN_16981; // @[rob.scala 124:83]
  wire  _GEN_19095 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12758 : _GEN_16982; // @[rob.scala 124:83]
  wire  _GEN_19096 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12759 : _GEN_16983; // @[rob.scala 124:83]
  wire  _GEN_19097 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12760 : _GEN_16984; // @[rob.scala 124:83]
  wire  _GEN_19098 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12761 : _GEN_16985; // @[rob.scala 124:83]
  wire  _GEN_19099 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12762 : _GEN_16986; // @[rob.scala 124:83]
  wire  _GEN_19100 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12763 : _GEN_16987; // @[rob.scala 124:83]
  wire  _GEN_19101 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12764 : _GEN_16988; // @[rob.scala 124:83]
  wire  _GEN_19102 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12765 : _GEN_16989; // @[rob.scala 124:83]
  wire  _GEN_19103 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12766 : _GEN_16990; // @[rob.scala 124:83]
  wire  _GEN_19104 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12767 : _GEN_16991; // @[rob.scala 124:83]
  wire  _GEN_19105 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12768 : _GEN_16992; // @[rob.scala 124:83]
  wire  _GEN_19106 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12769 : _GEN_16993; // @[rob.scala 124:83]
  wire  _GEN_19107 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12770 : _GEN_16994; // @[rob.scala 124:83]
  wire  _GEN_19108 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12771 : _GEN_16995; // @[rob.scala 124:83]
  wire  _GEN_19109 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12772 : _GEN_16996; // @[rob.scala 124:83]
  wire  _GEN_19110 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12773 : _GEN_16997; // @[rob.scala 124:83]
  wire  _GEN_19111 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12774 : _GEN_16998; // @[rob.scala 124:83]
  wire  _GEN_19112 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12775 : _GEN_16999; // @[rob.scala 124:83]
  wire  _GEN_19113 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12776 : _GEN_17000; // @[rob.scala 124:83]
  wire  _GEN_19114 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12777 : _GEN_17001; // @[rob.scala 124:83]
  wire  _GEN_19115 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12778 : _GEN_17002; // @[rob.scala 124:83]
  wire  _GEN_19116 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12779 : _GEN_17003; // @[rob.scala 124:83]
  wire  _GEN_19117 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12780 : _GEN_17004; // @[rob.scala 124:83]
  wire  _GEN_19118 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12781 : _GEN_17005; // @[rob.scala 124:83]
  wire  _GEN_19119 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12782 : _GEN_17006; // @[rob.scala 124:83]
  wire  _GEN_19120 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12783 : _GEN_17007; // @[rob.scala 124:83]
  wire  _GEN_19121 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12784 : _GEN_17008; // @[rob.scala 124:83]
  wire  _GEN_19122 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12785 : _GEN_17009; // @[rob.scala 124:83]
  wire  _GEN_19123 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12786 : _GEN_17010; // @[rob.scala 124:83]
  wire  _GEN_19124 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12787 : _GEN_17011; // @[rob.scala 124:83]
  wire  _GEN_19125 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12788 : _GEN_17012; // @[rob.scala 124:83]
  wire  _GEN_19126 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12789 : _GEN_17013; // @[rob.scala 124:83]
  wire  _GEN_19127 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12790 : _GEN_17014; // @[rob.scala 124:83]
  wire  _GEN_19128 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12791 : _GEN_17015; // @[rob.scala 124:83]
  wire  _GEN_19129 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12792 : _GEN_17016; // @[rob.scala 124:83]
  wire  _GEN_19130 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12793 : _GEN_17017; // @[rob.scala 124:83]
  wire  _GEN_19131 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12794 : _GEN_17018; // @[rob.scala 124:83]
  wire  _GEN_19132 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12795 : _GEN_17019; // @[rob.scala 124:83]
  wire  _GEN_19133 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12796 : _GEN_17020; // @[rob.scala 124:83]
  wire  _GEN_19134 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12797 : _GEN_17021; // @[rob.scala 124:83]
  wire  _GEN_19135 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12798 : _GEN_17022; // @[rob.scala 124:83]
  wire  _GEN_19136 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12799 : _GEN_17023; // @[rob.scala 124:83]
  wire  _GEN_19137 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12800 : _GEN_17025; // @[rob.scala 124:83]
  wire  _GEN_19138 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12801 : _GEN_17026; // @[rob.scala 124:83]
  wire  _GEN_19139 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12802 : _GEN_17027; // @[rob.scala 124:83]
  wire  _GEN_19140 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12803 : _GEN_17028; // @[rob.scala 124:83]
  wire  _GEN_19141 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12804 : _GEN_17029; // @[rob.scala 124:83]
  wire  _GEN_19142 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12805 : _GEN_17030; // @[rob.scala 124:83]
  wire  _GEN_19143 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12806 : _GEN_17031; // @[rob.scala 124:83]
  wire  _GEN_19144 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12807 : _GEN_17032; // @[rob.scala 124:83]
  wire  _GEN_19145 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12808 : _GEN_17033; // @[rob.scala 124:83]
  wire  _GEN_19146 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12809 : _GEN_17034; // @[rob.scala 124:83]
  wire  _GEN_19147 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12810 : _GEN_17035; // @[rob.scala 124:83]
  wire  _GEN_19148 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12811 : _GEN_17036; // @[rob.scala 124:83]
  wire  _GEN_19149 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12812 : _GEN_17037; // @[rob.scala 124:83]
  wire  _GEN_19150 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12813 : _GEN_17038; // @[rob.scala 124:83]
  wire  _GEN_19151 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12814 : _GEN_17039; // @[rob.scala 124:83]
  wire  _GEN_19152 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12815 : _GEN_17040; // @[rob.scala 124:83]
  wire  _GEN_19153 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12816 : _GEN_17041; // @[rob.scala 124:83]
  wire  _GEN_19154 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12817 : _GEN_17042; // @[rob.scala 124:83]
  wire  _GEN_19155 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12818 : _GEN_17043; // @[rob.scala 124:83]
  wire  _GEN_19156 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12819 : _GEN_17044; // @[rob.scala 124:83]
  wire  _GEN_19157 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12820 : _GEN_17045; // @[rob.scala 124:83]
  wire  _GEN_19158 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12821 : _GEN_17046; // @[rob.scala 124:83]
  wire  _GEN_19159 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12822 : _GEN_17047; // @[rob.scala 124:83]
  wire  _GEN_19160 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12823 : _GEN_17048; // @[rob.scala 124:83]
  wire  _GEN_19161 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12824 : _GEN_17049; // @[rob.scala 124:83]
  wire  _GEN_19162 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12825 : _GEN_17050; // @[rob.scala 124:83]
  wire  _GEN_19163 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12826 : _GEN_17051; // @[rob.scala 124:83]
  wire  _GEN_19164 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12827 : _GEN_17052; // @[rob.scala 124:83]
  wire  _GEN_19165 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12828 : _GEN_17053; // @[rob.scala 124:83]
  wire  _GEN_19166 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12829 : _GEN_17054; // @[rob.scala 124:83]
  wire  _GEN_19167 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12830 : _GEN_17055; // @[rob.scala 124:83]
  wire  _GEN_19168 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12831 : _GEN_17056; // @[rob.scala 124:83]
  wire  _GEN_19169 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12832 : _GEN_17057; // @[rob.scala 124:83]
  wire  _GEN_19170 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12833 : _GEN_17058; // @[rob.scala 124:83]
  wire  _GEN_19171 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12834 : _GEN_17059; // @[rob.scala 124:83]
  wire  _GEN_19172 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12835 : _GEN_17060; // @[rob.scala 124:83]
  wire  _GEN_19173 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12836 : _GEN_17061; // @[rob.scala 124:83]
  wire  _GEN_19174 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12837 : _GEN_17062; // @[rob.scala 124:83]
  wire  _GEN_19175 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12838 : _GEN_17063; // @[rob.scala 124:83]
  wire  _GEN_19176 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12839 : _GEN_17064; // @[rob.scala 124:83]
  wire  _GEN_19177 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12840 : _GEN_17065; // @[rob.scala 124:83]
  wire  _GEN_19178 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12841 : _GEN_17066; // @[rob.scala 124:83]
  wire  _GEN_19179 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12842 : _GEN_17067; // @[rob.scala 124:83]
  wire  _GEN_19180 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12843 : _GEN_17068; // @[rob.scala 124:83]
  wire  _GEN_19181 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12844 : _GEN_17069; // @[rob.scala 124:83]
  wire  _GEN_19182 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12845 : _GEN_17070; // @[rob.scala 124:83]
  wire  _GEN_19183 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12846 : _GEN_17071; // @[rob.scala 124:83]
  wire  _GEN_19184 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12847 : _GEN_17072; // @[rob.scala 124:83]
  wire  _GEN_19185 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12848 : _GEN_17073; // @[rob.scala 124:83]
  wire  _GEN_19186 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12849 : _GEN_17074; // @[rob.scala 124:83]
  wire  _GEN_19187 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12850 : _GEN_17075; // @[rob.scala 124:83]
  wire  _GEN_19188 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12851 : _GEN_17076; // @[rob.scala 124:83]
  wire  _GEN_19189 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12852 : _GEN_17077; // @[rob.scala 124:83]
  wire  _GEN_19190 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12853 : _GEN_17078; // @[rob.scala 124:83]
  wire  _GEN_19191 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12854 : _GEN_17079; // @[rob.scala 124:83]
  wire  _GEN_19192 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12855 : _GEN_17080; // @[rob.scala 124:83]
  wire  _GEN_19193 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12856 : _GEN_17081; // @[rob.scala 124:83]
  wire  _GEN_19194 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12857 : _GEN_17082; // @[rob.scala 124:83]
  wire  _GEN_19195 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12858 : _GEN_17083; // @[rob.scala 124:83]
  wire  _GEN_19196 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12859 : _GEN_17084; // @[rob.scala 124:83]
  wire  _GEN_19197 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12860 : _GEN_17085; // @[rob.scala 124:83]
  wire  _GEN_19198 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12861 : _GEN_17086; // @[rob.scala 124:83]
  wire  _GEN_19199 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12862 : _GEN_17087; // @[rob.scala 124:83]
  wire  _GEN_19200 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _GEN_12863 : _GEN_17088; // @[rob.scala 124:83]
  wire [6:0] _GEN_19201 = io_i_rob_allocation_reqs_0_valid & io_i_rob_allocation_reqs_1_valid ? _is_full_T_1 :
    _GEN_17024; // @[rob.scala 124:83 132:22]
  wire  _GEN_42065 = 6'h0 == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19202 = 6'h0 == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19073; // @[rob.scala 142:{53,53}]
  wire  _GEN_42066 = 6'h1 == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19203 = 6'h1 == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19074; // @[rob.scala 142:{53,53}]
  wire  _GEN_42067 = 6'h2 == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19204 = 6'h2 == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19075; // @[rob.scala 142:{53,53}]
  wire  _GEN_42068 = 6'h3 == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19205 = 6'h3 == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19076; // @[rob.scala 142:{53,53}]
  wire  _GEN_42069 = 6'h4 == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19206 = 6'h4 == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19077; // @[rob.scala 142:{53,53}]
  wire  _GEN_42070 = 6'h5 == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19207 = 6'h5 == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19078; // @[rob.scala 142:{53,53}]
  wire  _GEN_42071 = 6'h6 == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19208 = 6'h6 == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19079; // @[rob.scala 142:{53,53}]
  wire  _GEN_42072 = 6'h7 == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19209 = 6'h7 == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19080; // @[rob.scala 142:{53,53}]
  wire  _GEN_42073 = 6'h8 == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19210 = 6'h8 == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19081; // @[rob.scala 142:{53,53}]
  wire  _GEN_42074 = 6'h9 == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19211 = 6'h9 == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19082; // @[rob.scala 142:{53,53}]
  wire  _GEN_42075 = 6'ha == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19212 = 6'ha == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19083; // @[rob.scala 142:{53,53}]
  wire  _GEN_42076 = 6'hb == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19213 = 6'hb == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19084; // @[rob.scala 142:{53,53}]
  wire  _GEN_42077 = 6'hc == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19214 = 6'hc == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19085; // @[rob.scala 142:{53,53}]
  wire  _GEN_42078 = 6'hd == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19215 = 6'hd == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19086; // @[rob.scala 142:{53,53}]
  wire  _GEN_42079 = 6'he == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19216 = 6'he == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19087; // @[rob.scala 142:{53,53}]
  wire  _GEN_42080 = 6'hf == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19217 = 6'hf == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19088; // @[rob.scala 142:{53,53}]
  wire  _GEN_42081 = 6'h10 == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19218 = 6'h10 == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19089; // @[rob.scala 142:{53,53}]
  wire  _GEN_42082 = 6'h11 == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19219 = 6'h11 == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19090; // @[rob.scala 142:{53,53}]
  wire  _GEN_42083 = 6'h12 == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19220 = 6'h12 == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19091; // @[rob.scala 142:{53,53}]
  wire  _GEN_42084 = 6'h13 == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19221 = 6'h13 == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19092; // @[rob.scala 142:{53,53}]
  wire  _GEN_42085 = 6'h14 == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19222 = 6'h14 == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19093; // @[rob.scala 142:{53,53}]
  wire  _GEN_42086 = 6'h15 == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19223 = 6'h15 == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19094; // @[rob.scala 142:{53,53}]
  wire  _GEN_42087 = 6'h16 == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19224 = 6'h16 == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19095; // @[rob.scala 142:{53,53}]
  wire  _GEN_42088 = 6'h17 == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19225 = 6'h17 == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19096; // @[rob.scala 142:{53,53}]
  wire  _GEN_42089 = 6'h18 == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19226 = 6'h18 == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19097; // @[rob.scala 142:{53,53}]
  wire  _GEN_42090 = 6'h19 == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19227 = 6'h19 == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19098; // @[rob.scala 142:{53,53}]
  wire  _GEN_42091 = 6'h1a == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19228 = 6'h1a == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19099; // @[rob.scala 142:{53,53}]
  wire  _GEN_42092 = 6'h1b == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19229 = 6'h1b == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19100; // @[rob.scala 142:{53,53}]
  wire  _GEN_42093 = 6'h1c == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19230 = 6'h1c == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19101; // @[rob.scala 142:{53,53}]
  wire  _GEN_42094 = 6'h1d == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19231 = 6'h1d == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19102; // @[rob.scala 142:{53,53}]
  wire  _GEN_42095 = 6'h1e == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19232 = 6'h1e == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19103; // @[rob.scala 142:{53,53}]
  wire  _GEN_42096 = 6'h1f == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19233 = 6'h1f == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19104; // @[rob.scala 142:{53,53}]
  wire  _GEN_42097 = 6'h20 == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19234 = 6'h20 == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19105; // @[rob.scala 142:{53,53}]
  wire  _GEN_42098 = 6'h21 == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19235 = 6'h21 == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19106; // @[rob.scala 142:{53,53}]
  wire  _GEN_42099 = 6'h22 == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19236 = 6'h22 == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19107; // @[rob.scala 142:{53,53}]
  wire  _GEN_42100 = 6'h23 == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19237 = 6'h23 == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19108; // @[rob.scala 142:{53,53}]
  wire  _GEN_42101 = 6'h24 == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19238 = 6'h24 == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19109; // @[rob.scala 142:{53,53}]
  wire  _GEN_42102 = 6'h25 == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19239 = 6'h25 == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19110; // @[rob.scala 142:{53,53}]
  wire  _GEN_42103 = 6'h26 == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19240 = 6'h26 == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19111; // @[rob.scala 142:{53,53}]
  wire  _GEN_42104 = 6'h27 == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19241 = 6'h27 == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19112; // @[rob.scala 142:{53,53}]
  wire  _GEN_42105 = 6'h28 == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19242 = 6'h28 == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19113; // @[rob.scala 142:{53,53}]
  wire  _GEN_42106 = 6'h29 == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19243 = 6'h29 == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19114; // @[rob.scala 142:{53,53}]
  wire  _GEN_42107 = 6'h2a == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19244 = 6'h2a == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19115; // @[rob.scala 142:{53,53}]
  wire  _GEN_42108 = 6'h2b == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19245 = 6'h2b == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19116; // @[rob.scala 142:{53,53}]
  wire  _GEN_42109 = 6'h2c == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19246 = 6'h2c == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19117; // @[rob.scala 142:{53,53}]
  wire  _GEN_42110 = 6'h2d == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19247 = 6'h2d == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19118; // @[rob.scala 142:{53,53}]
  wire  _GEN_42111 = 6'h2e == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19248 = 6'h2e == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19119; // @[rob.scala 142:{53,53}]
  wire  _GEN_42112 = 6'h2f == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19249 = 6'h2f == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19120; // @[rob.scala 142:{53,53}]
  wire  _GEN_42113 = 6'h30 == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19250 = 6'h30 == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19121; // @[rob.scala 142:{53,53}]
  wire  _GEN_42114 = 6'h31 == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19251 = 6'h31 == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19122; // @[rob.scala 142:{53,53}]
  wire  _GEN_42115 = 6'h32 == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19252 = 6'h32 == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19123; // @[rob.scala 142:{53,53}]
  wire  _GEN_42116 = 6'h33 == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19253 = 6'h33 == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19124; // @[rob.scala 142:{53,53}]
  wire  _GEN_42117 = 6'h34 == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19254 = 6'h34 == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19125; // @[rob.scala 142:{53,53}]
  wire  _GEN_42118 = 6'h35 == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19255 = 6'h35 == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19126; // @[rob.scala 142:{53,53}]
  wire  _GEN_42119 = 6'h36 == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19256 = 6'h36 == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19127; // @[rob.scala 142:{53,53}]
  wire  _GEN_42120 = 6'h37 == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19257 = 6'h37 == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19128; // @[rob.scala 142:{53,53}]
  wire  _GEN_42121 = 6'h38 == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19258 = 6'h38 == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19129; // @[rob.scala 142:{53,53}]
  wire  _GEN_42122 = 6'h39 == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19259 = 6'h39 == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19130; // @[rob.scala 142:{53,53}]
  wire  _GEN_42123 = 6'h3a == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19260 = 6'h3a == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19131; // @[rob.scala 142:{53,53}]
  wire  _GEN_42124 = 6'h3b == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19261 = 6'h3b == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19132; // @[rob.scala 142:{53,53}]
  wire  _GEN_42125 = 6'h3c == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19262 = 6'h3c == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19133; // @[rob.scala 142:{53,53}]
  wire  _GEN_42126 = 6'h3d == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19263 = 6'h3d == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19134; // @[rob.scala 142:{53,53}]
  wire  _GEN_42127 = 6'h3e == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19264 = 6'h3e == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19135; // @[rob.scala 142:{53,53}]
  wire  _GEN_42128 = 6'h3f == io_i_ex_res_packs_0_uop_rob_idx[5:0]; // @[rob.scala 142:{53,53}]
  wire  _GEN_19265 = 6'h3f == io_i_ex_res_packs_0_uop_rob_idx[5:0] | _GEN_19136; // @[rob.scala 142:{53,53}]
  wire [31:0] _GEN_19330 = 6'h0 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17153; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19331 = 6'h1 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17154; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19332 = 6'h2 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17155; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19333 = 6'h3 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17156; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19334 = 6'h4 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17157; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19335 = 6'h5 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17158; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19336 = 6'h6 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17159; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19337 = 6'h7 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17160; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19338 = 6'h8 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17161; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19339 = 6'h9 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17162; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19340 = 6'ha == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17163; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19341 = 6'hb == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17164; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19342 = 6'hc == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17165; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19343 = 6'hd == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17166; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19344 = 6'he == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17167; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19345 = 6'hf == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17168; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19346 = 6'h10 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17169; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19347 = 6'h11 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17170; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19348 = 6'h12 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17171; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19349 = 6'h13 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17172; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19350 = 6'h14 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17173; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19351 = 6'h15 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17174; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19352 = 6'h16 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17175; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19353 = 6'h17 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17176; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19354 = 6'h18 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17177; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19355 = 6'h19 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17178; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19356 = 6'h1a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17179; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19357 = 6'h1b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17180; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19358 = 6'h1c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17181; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19359 = 6'h1d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17182; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19360 = 6'h1e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17183; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19361 = 6'h1f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17184; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19362 = 6'h20 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17185; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19363 = 6'h21 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17186; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19364 = 6'h22 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17187; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19365 = 6'h23 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17188; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19366 = 6'h24 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17189; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19367 = 6'h25 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17190; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19368 = 6'h26 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17191; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19369 = 6'h27 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17192; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19370 = 6'h28 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17193; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19371 = 6'h29 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17194; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19372 = 6'h2a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17195; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19373 = 6'h2b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17196; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19374 = 6'h2c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17197; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19375 = 6'h2d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17198; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19376 = 6'h2e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17199; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19377 = 6'h2f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17200; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19378 = 6'h30 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17201; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19379 = 6'h31 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17202; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19380 = 6'h32 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17203; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19381 = 6'h33 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17204; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19382 = 6'h34 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17205; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19383 = 6'h35 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17206; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19384 = 6'h36 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17207; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19385 = 6'h37 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17208; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19386 = 6'h38 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17209; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19387 = 6'h39 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17210; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19388 = 6'h3a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17211; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19389 = 6'h3b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17212; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19390 = 6'h3c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17213; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19391 = 6'h3d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17214; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19392 = 6'h3e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17215; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19393 = 6'h3f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_17216; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19394 = 6'h0 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17217; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19395 = 6'h1 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17218; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19396 = 6'h2 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17219; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19397 = 6'h3 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17220; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19398 = 6'h4 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17221; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19399 = 6'h5 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17222; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19400 = 6'h6 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17223; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19401 = 6'h7 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17224; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19402 = 6'h8 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17225; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19403 = 6'h9 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17226; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19404 = 6'ha == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17227; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19405 = 6'hb == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17228; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19406 = 6'hc == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17229; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19407 = 6'hd == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17230; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19408 = 6'he == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17231; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19409 = 6'hf == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17232; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19410 = 6'h10 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17233; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19411 = 6'h11 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17234; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19412 = 6'h12 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17235; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19413 = 6'h13 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17236; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19414 = 6'h14 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17237; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19415 = 6'h15 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17238; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19416 = 6'h16 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17239; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19417 = 6'h17 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17240; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19418 = 6'h18 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17241; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19419 = 6'h19 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17242; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19420 = 6'h1a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17243; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19421 = 6'h1b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17244; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19422 = 6'h1c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17245; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19423 = 6'h1d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17246; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19424 = 6'h1e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17247; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19425 = 6'h1f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17248; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19426 = 6'h20 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17249; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19427 = 6'h21 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17250; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19428 = 6'h22 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17251; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19429 = 6'h23 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17252; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19430 = 6'h24 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17253; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19431 = 6'h25 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17254; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19432 = 6'h26 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17255; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19433 = 6'h27 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17256; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19434 = 6'h28 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17257; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19435 = 6'h29 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17258; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19436 = 6'h2a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17259; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19437 = 6'h2b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17260; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19438 = 6'h2c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17261; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19439 = 6'h2d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17262; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19440 = 6'h2e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17263; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19441 = 6'h2f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17264; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19442 = 6'h30 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17265; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19443 = 6'h31 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17266; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19444 = 6'h32 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17267; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19445 = 6'h33 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17268; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19446 = 6'h34 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17269; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19447 = 6'h35 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17270; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19448 = 6'h36 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17271; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19449 = 6'h37 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17272; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19450 = 6'h38 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17273; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19451 = 6'h39 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17274; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19452 = 6'h3a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17275; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19453 = 6'h3b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17276; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19454 = 6'h3c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17277; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19455 = 6'h3d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17278; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19456 = 6'h3e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17279; // @[rob.scala 143:{51,51}]
  wire [31:0] _GEN_19457 = 6'h3f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_17280; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19458 = 6'h0 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17281; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19459 = 6'h1 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17282; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19460 = 6'h2 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17283; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19461 = 6'h3 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17284; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19462 = 6'h4 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17285; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19463 = 6'h5 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17286; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19464 = 6'h6 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17287; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19465 = 6'h7 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17288; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19466 = 6'h8 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17289; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19467 = 6'h9 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17290; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19468 = 6'ha == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17291; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19469 = 6'hb == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17292; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19470 = 6'hc == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17293; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19471 = 6'hd == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17294; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19472 = 6'he == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17295; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19473 = 6'hf == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17296; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19474 = 6'h10 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17297
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19475 = 6'h11 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17298
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19476 = 6'h12 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17299
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19477 = 6'h13 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17300
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19478 = 6'h14 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17301
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19479 = 6'h15 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17302
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19480 = 6'h16 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17303
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19481 = 6'h17 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17304
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19482 = 6'h18 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17305
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19483 = 6'h19 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17306
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19484 = 6'h1a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17307
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19485 = 6'h1b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17308
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19486 = 6'h1c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17309
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19487 = 6'h1d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17310
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19488 = 6'h1e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17311
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19489 = 6'h1f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17312
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19490 = 6'h20 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17313
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19491 = 6'h21 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17314
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19492 = 6'h22 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17315
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19493 = 6'h23 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17316
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19494 = 6'h24 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17317
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19495 = 6'h25 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17318
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19496 = 6'h26 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17319
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19497 = 6'h27 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17320
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19498 = 6'h28 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17321
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19499 = 6'h29 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17322
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19500 = 6'h2a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17323
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19501 = 6'h2b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17324
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19502 = 6'h2c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17325
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19503 = 6'h2d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17326
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19504 = 6'h2e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17327
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19505 = 6'h2f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17328
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19506 = 6'h30 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17329
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19507 = 6'h31 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17330
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19508 = 6'h32 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17331
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19509 = 6'h33 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17332
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19510 = 6'h34 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17333
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19511 = 6'h35 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17334
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19512 = 6'h36 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17335
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19513 = 6'h37 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17336
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19514 = 6'h38 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17337
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19515 = 6'h39 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17338
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19516 = 6'h3a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17339
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19517 = 6'h3b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17340
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19518 = 6'h3c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17341
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19519 = 6'h3d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17342
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19520 = 6'h3e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17343
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19521 = 6'h3f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_17344
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19842 = 6'h0 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17665; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19843 = 6'h1 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17666; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19844 = 6'h2 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17667; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19845 = 6'h3 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17668; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19846 = 6'h4 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17669; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19847 = 6'h5 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17670; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19848 = 6'h6 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17671; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19849 = 6'h7 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17672; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19850 = 6'h8 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17673; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19851 = 6'h9 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17674; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19852 = 6'ha == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17675; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19853 = 6'hb == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17676; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19854 = 6'hc == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17677; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19855 = 6'hd == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17678; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19856 = 6'he == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17679; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19857 = 6'hf == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17680; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19858 = 6'h10 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17681; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19859 = 6'h11 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17682; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19860 = 6'h12 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17683; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19861 = 6'h13 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17684; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19862 = 6'h14 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17685; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19863 = 6'h15 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17686; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19864 = 6'h16 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17687; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19865 = 6'h17 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17688; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19866 = 6'h18 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17689; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19867 = 6'h19 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17690; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19868 = 6'h1a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17691; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19869 = 6'h1b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17692; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19870 = 6'h1c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17693; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19871 = 6'h1d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17694; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19872 = 6'h1e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17695; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19873 = 6'h1f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17696; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19874 = 6'h20 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17697; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19875 = 6'h21 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17698; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19876 = 6'h22 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17699; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19877 = 6'h23 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17700; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19878 = 6'h24 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17701; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19879 = 6'h25 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17702; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19880 = 6'h26 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17703; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19881 = 6'h27 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17704; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19882 = 6'h28 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17705; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19883 = 6'h29 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17706; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19884 = 6'h2a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17707; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19885 = 6'h2b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17708; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19886 = 6'h2c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17709; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19887 = 6'h2d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17710; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19888 = 6'h2e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17711; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19889 = 6'h2f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17712; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19890 = 6'h30 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17713; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19891 = 6'h31 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17714; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19892 = 6'h32 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17715; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19893 = 6'h33 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17716; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19894 = 6'h34 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17717; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19895 = 6'h35 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17718; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19896 = 6'h36 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17719; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19897 = 6'h37 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17720; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19898 = 6'h38 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17721; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19899 = 6'h39 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17722; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19900 = 6'h3a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17723; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19901 = 6'h3b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17724; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19902 = 6'h3c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17725; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19903 = 6'h3d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17726; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19904 = 6'h3e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17727; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19905 = 6'h3f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_17728; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19906 = 6'h0 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17729; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19907 = 6'h1 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17730; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19908 = 6'h2 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17731; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19909 = 6'h3 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17732; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19910 = 6'h4 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17733; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19911 = 6'h5 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17734; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19912 = 6'h6 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17735; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19913 = 6'h7 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17736; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19914 = 6'h8 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17737; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19915 = 6'h9 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17738; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19916 = 6'ha == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17739; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19917 = 6'hb == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17740; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19918 = 6'hc == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17741; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19919 = 6'hd == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17742; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19920 = 6'he == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17743; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19921 = 6'hf == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17744; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19922 = 6'h10 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17745
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19923 = 6'h11 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17746
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19924 = 6'h12 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17747
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19925 = 6'h13 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17748
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19926 = 6'h14 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17749
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19927 = 6'h15 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17750
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19928 = 6'h16 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17751
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19929 = 6'h17 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17752
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19930 = 6'h18 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17753
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19931 = 6'h19 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17754
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19932 = 6'h1a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17755
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19933 = 6'h1b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17756
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19934 = 6'h1c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17757
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19935 = 6'h1d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17758
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19936 = 6'h1e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17759
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19937 = 6'h1f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17760
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19938 = 6'h20 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17761
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19939 = 6'h21 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17762
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19940 = 6'h22 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17763
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19941 = 6'h23 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17764
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19942 = 6'h24 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17765
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19943 = 6'h25 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17766
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19944 = 6'h26 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17767
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19945 = 6'h27 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17768
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19946 = 6'h28 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17769
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19947 = 6'h29 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17770
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19948 = 6'h2a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17771
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19949 = 6'h2b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17772
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19950 = 6'h2c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17773
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19951 = 6'h2d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17774
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19952 = 6'h2e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17775
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19953 = 6'h2f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17776
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19954 = 6'h30 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17777
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19955 = 6'h31 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17778
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19956 = 6'h32 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17779
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19957 = 6'h33 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17780
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19958 = 6'h34 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17781
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19959 = 6'h35 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17782
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19960 = 6'h36 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17783
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19961 = 6'h37 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17784
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19962 = 6'h38 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17785
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19963 = 6'h39 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17786
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19964 = 6'h3a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17787
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19965 = 6'h3b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17788
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19966 = 6'h3c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17789
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19967 = 6'h3d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17790
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19968 = 6'h3e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17791
    ; // @[rob.scala 143:{51,51}]
  wire [6:0] _GEN_19969 = 6'h3f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_17792
    ; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_19970 = 6'h0 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17793; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_19971 = 6'h1 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17794; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_19972 = 6'h2 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17795; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_19973 = 6'h3 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17796; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_19974 = 6'h4 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17797; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_19975 = 6'h5 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17798; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_19976 = 6'h6 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17799; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_19977 = 6'h7 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17800; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_19978 = 6'h8 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17801; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_19979 = 6'h9 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17802; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_19980 = 6'ha == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17803; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_19981 = 6'hb == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17804; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_19982 = 6'hc == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17805; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_19983 = 6'hd == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17806; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_19984 = 6'he == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17807; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_19985 = 6'hf == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17808; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_19986 = 6'h10 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17809; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_19987 = 6'h11 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17810; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_19988 = 6'h12 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17811; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_19989 = 6'h13 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17812; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_19990 = 6'h14 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17813; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_19991 = 6'h15 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17814; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_19992 = 6'h16 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17815; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_19993 = 6'h17 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17816; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_19994 = 6'h18 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17817; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_19995 = 6'h19 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17818; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_19996 = 6'h1a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17819; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_19997 = 6'h1b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17820; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_19998 = 6'h1c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17821; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_19999 = 6'h1d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17822; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_20000 = 6'h1e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17823; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_20001 = 6'h1f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17824; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_20002 = 6'h20 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17825; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_20003 = 6'h21 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17826; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_20004 = 6'h22 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17827; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_20005 = 6'h23 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17828; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_20006 = 6'h24 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17829; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_20007 = 6'h25 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17830; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_20008 = 6'h26 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17831; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_20009 = 6'h27 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17832; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_20010 = 6'h28 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17833; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_20011 = 6'h29 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17834; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_20012 = 6'h2a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17835; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_20013 = 6'h2b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17836; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_20014 = 6'h2c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17837; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_20015 = 6'h2d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17838; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_20016 = 6'h2e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17839; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_20017 = 6'h2f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17840; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_20018 = 6'h30 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17841; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_20019 = 6'h31 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17842; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_20020 = 6'h32 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17843; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_20021 = 6'h33 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17844; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_20022 = 6'h34 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17845; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_20023 = 6'h35 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17846; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_20024 = 6'h36 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17847; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_20025 = 6'h37 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17848; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_20026 = 6'h38 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17849; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_20027 = 6'h39 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17850; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_20028 = 6'h3a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17851; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_20029 = 6'h3b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17852; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_20030 = 6'h3c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17853; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_20031 = 6'h3d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17854; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_20032 = 6'h3e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17855; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_20033 = 6'h3f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_17856; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20674 = 6'h0 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value : _GEN_18497
    ; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20675 = 6'h1 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value : _GEN_18498
    ; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20676 = 6'h2 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value : _GEN_18499
    ; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20677 = 6'h3 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value : _GEN_18500
    ; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20678 = 6'h4 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value : _GEN_18501
    ; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20679 = 6'h5 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value : _GEN_18502
    ; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20680 = 6'h6 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value : _GEN_18503
    ; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20681 = 6'h7 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value : _GEN_18504
    ; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20682 = 6'h8 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value : _GEN_18505
    ; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20683 = 6'h9 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value : _GEN_18506
    ; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20684 = 6'ha == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value : _GEN_18507
    ; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20685 = 6'hb == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value : _GEN_18508
    ; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20686 = 6'hc == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value : _GEN_18509
    ; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20687 = 6'hd == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value : _GEN_18510
    ; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20688 = 6'he == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value : _GEN_18511
    ; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20689 = 6'hf == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value : _GEN_18512
    ; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20690 = 6'h10 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18513; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20691 = 6'h11 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18514; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20692 = 6'h12 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18515; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20693 = 6'h13 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18516; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20694 = 6'h14 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18517; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20695 = 6'h15 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18518; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20696 = 6'h16 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18519; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20697 = 6'h17 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18520; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20698 = 6'h18 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18521; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20699 = 6'h19 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18522; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20700 = 6'h1a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18523; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20701 = 6'h1b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18524; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20702 = 6'h1c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18525; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20703 = 6'h1d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18526; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20704 = 6'h1e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18527; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20705 = 6'h1f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18528; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20706 = 6'h20 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18529; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20707 = 6'h21 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18530; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20708 = 6'h22 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18531; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20709 = 6'h23 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18532; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20710 = 6'h24 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18533; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20711 = 6'h25 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18534; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20712 = 6'h26 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18535; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20713 = 6'h27 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18536; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20714 = 6'h28 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18537; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20715 = 6'h29 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18538; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20716 = 6'h2a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18539; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20717 = 6'h2b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18540; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20718 = 6'h2c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18541; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20719 = 6'h2d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18542; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20720 = 6'h2e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18543; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20721 = 6'h2f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18544; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20722 = 6'h30 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18545; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20723 = 6'h31 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18546; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20724 = 6'h32 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18547; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20725 = 6'h33 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18548; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20726 = 6'h34 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18549; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20727 = 6'h35 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18550; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20728 = 6'h36 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18551; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20729 = 6'h37 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18552; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20730 = 6'h38 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18553; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20731 = 6'h39 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18554; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20732 = 6'h3a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18555; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20733 = 6'h3b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18556; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20734 = 6'h3c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18557; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20735 = 6'h3d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18558; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20736 = 6'h3e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18559; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20737 = 6'h3f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_18560; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20738 = 6'h0 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18561; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20739 = 6'h1 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18562; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20740 = 6'h2 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18563; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20741 = 6'h3 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18564; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20742 = 6'h4 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18565; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20743 = 6'h5 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18566; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20744 = 6'h6 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18567; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20745 = 6'h7 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18568; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20746 = 6'h8 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18569; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20747 = 6'h9 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18570; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20748 = 6'ha == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18571; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20749 = 6'hb == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18572; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20750 = 6'hc == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18573; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20751 = 6'hd == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18574; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20752 = 6'he == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18575; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20753 = 6'hf == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18576; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20754 = 6'h10 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18577; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20755 = 6'h11 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18578; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20756 = 6'h12 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18579; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20757 = 6'h13 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18580; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20758 = 6'h14 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18581; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20759 = 6'h15 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18582; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20760 = 6'h16 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18583; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20761 = 6'h17 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18584; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20762 = 6'h18 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18585; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20763 = 6'h19 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18586; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20764 = 6'h1a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18587; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20765 = 6'h1b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18588; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20766 = 6'h1c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18589; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20767 = 6'h1d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18590; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20768 = 6'h1e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18591; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20769 = 6'h1f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18592; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20770 = 6'h20 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18593; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20771 = 6'h21 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18594; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20772 = 6'h22 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18595; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20773 = 6'h23 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18596; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20774 = 6'h24 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18597; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20775 = 6'h25 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18598; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20776 = 6'h26 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18599; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20777 = 6'h27 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18600; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20778 = 6'h28 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18601; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20779 = 6'h29 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18602; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20780 = 6'h2a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18603; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20781 = 6'h2b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18604; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20782 = 6'h2c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18605; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20783 = 6'h2d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18606; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20784 = 6'h2e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18607; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20785 = 6'h2f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18608; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20786 = 6'h30 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18609; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20787 = 6'h31 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18610; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20788 = 6'h32 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18611; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20789 = 6'h33 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18612; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20790 = 6'h34 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18613; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20791 = 6'h35 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18614; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20792 = 6'h36 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18615; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20793 = 6'h37 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18616; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20794 = 6'h38 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18617; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20795 = 6'h39 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18618; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20796 = 6'h3a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18619; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20797 = 6'h3b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18620; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20798 = 6'h3c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18621; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20799 = 6'h3d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18622; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20800 = 6'h3e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18623; // @[rob.scala 143:{51,51}]
  wire [63:0] _GEN_20801 = 6'h3f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_18624; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21058 = 6'h0 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18881; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21059 = 6'h1 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18882; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21060 = 6'h2 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18883; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21061 = 6'h3 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18884; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21062 = 6'h4 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18885; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21063 = 6'h5 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18886; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21064 = 6'h6 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18887; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21065 = 6'h7 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18888; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21066 = 6'h8 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18889; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21067 = 6'h9 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18890; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21068 = 6'ha == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18891; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21069 = 6'hb == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18892; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21070 = 6'hc == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18893; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21071 = 6'hd == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18894; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21072 = 6'he == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18895; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21073 = 6'hf == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18896; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21074 = 6'h10 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18897; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21075 = 6'h11 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18898; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21076 = 6'h12 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18899; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21077 = 6'h13 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18900; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21078 = 6'h14 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18901; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21079 = 6'h15 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18902; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21080 = 6'h16 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18903; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21081 = 6'h17 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18904; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21082 = 6'h18 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18905; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21083 = 6'h19 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18906; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21084 = 6'h1a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18907; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21085 = 6'h1b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18908; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21086 = 6'h1c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18909; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21087 = 6'h1d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18910; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21088 = 6'h1e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18911; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21089 = 6'h1f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18912; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21090 = 6'h20 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18913; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21091 = 6'h21 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18914; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21092 = 6'h22 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18915; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21093 = 6'h23 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18916; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21094 = 6'h24 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18917; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21095 = 6'h25 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18918; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21096 = 6'h26 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18919; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21097 = 6'h27 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18920; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21098 = 6'h28 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18921; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21099 = 6'h29 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18922; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21100 = 6'h2a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18923; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21101 = 6'h2b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18924; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21102 = 6'h2c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18925; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21103 = 6'h2d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18926; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21104 = 6'h2e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18927; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21105 = 6'h2f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18928; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21106 = 6'h30 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18929; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21107 = 6'h31 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18930; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21108 = 6'h32 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18931; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21109 = 6'h33 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18932; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21110 = 6'h34 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18933; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21111 = 6'h35 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18934; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21112 = 6'h36 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18935; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21113 = 6'h37 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18936; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21114 = 6'h38 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18937; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21115 = 6'h39 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18938; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21116 = 6'h3a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18939; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21117 = 6'h3b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18940; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21118 = 6'h3c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18941; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21119 = 6'h3d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18942; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21120 = 6'h3e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18943; // @[rob.scala 143:{51,51}]
  wire [4:0] _GEN_21121 = 6'h3f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_18944; // @[rob.scala 143:{51,51}]
  wire  _GEN_21314 = _GEN_42065 | _GEN_19137; // @[rob.scala 145:{52,52}]
  wire  _GEN_21315 = _GEN_42066 | _GEN_19138; // @[rob.scala 145:{52,52}]
  wire  _GEN_21316 = _GEN_42067 | _GEN_19139; // @[rob.scala 145:{52,52}]
  wire  _GEN_21317 = _GEN_42068 | _GEN_19140; // @[rob.scala 145:{52,52}]
  wire  _GEN_21318 = _GEN_42069 | _GEN_19141; // @[rob.scala 145:{52,52}]
  wire  _GEN_21319 = _GEN_42070 | _GEN_19142; // @[rob.scala 145:{52,52}]
  wire  _GEN_21320 = _GEN_42071 | _GEN_19143; // @[rob.scala 145:{52,52}]
  wire  _GEN_21321 = _GEN_42072 | _GEN_19144; // @[rob.scala 145:{52,52}]
  wire  _GEN_21322 = _GEN_42073 | _GEN_19145; // @[rob.scala 145:{52,52}]
  wire  _GEN_21323 = _GEN_42074 | _GEN_19146; // @[rob.scala 145:{52,52}]
  wire  _GEN_21324 = _GEN_42075 | _GEN_19147; // @[rob.scala 145:{52,52}]
  wire  _GEN_21325 = _GEN_42076 | _GEN_19148; // @[rob.scala 145:{52,52}]
  wire  _GEN_21326 = _GEN_42077 | _GEN_19149; // @[rob.scala 145:{52,52}]
  wire  _GEN_21327 = _GEN_42078 | _GEN_19150; // @[rob.scala 145:{52,52}]
  wire  _GEN_21328 = _GEN_42079 | _GEN_19151; // @[rob.scala 145:{52,52}]
  wire  _GEN_21329 = _GEN_42080 | _GEN_19152; // @[rob.scala 145:{52,52}]
  wire  _GEN_21330 = _GEN_42081 | _GEN_19153; // @[rob.scala 145:{52,52}]
  wire  _GEN_21331 = _GEN_42082 | _GEN_19154; // @[rob.scala 145:{52,52}]
  wire  _GEN_21332 = _GEN_42083 | _GEN_19155; // @[rob.scala 145:{52,52}]
  wire  _GEN_21333 = _GEN_42084 | _GEN_19156; // @[rob.scala 145:{52,52}]
  wire  _GEN_21334 = _GEN_42085 | _GEN_19157; // @[rob.scala 145:{52,52}]
  wire  _GEN_21335 = _GEN_42086 | _GEN_19158; // @[rob.scala 145:{52,52}]
  wire  _GEN_21336 = _GEN_42087 | _GEN_19159; // @[rob.scala 145:{52,52}]
  wire  _GEN_21337 = _GEN_42088 | _GEN_19160; // @[rob.scala 145:{52,52}]
  wire  _GEN_21338 = _GEN_42089 | _GEN_19161; // @[rob.scala 145:{52,52}]
  wire  _GEN_21339 = _GEN_42090 | _GEN_19162; // @[rob.scala 145:{52,52}]
  wire  _GEN_21340 = _GEN_42091 | _GEN_19163; // @[rob.scala 145:{52,52}]
  wire  _GEN_21341 = _GEN_42092 | _GEN_19164; // @[rob.scala 145:{52,52}]
  wire  _GEN_21342 = _GEN_42093 | _GEN_19165; // @[rob.scala 145:{52,52}]
  wire  _GEN_21343 = _GEN_42094 | _GEN_19166; // @[rob.scala 145:{52,52}]
  wire  _GEN_21344 = _GEN_42095 | _GEN_19167; // @[rob.scala 145:{52,52}]
  wire  _GEN_21345 = _GEN_42096 | _GEN_19168; // @[rob.scala 145:{52,52}]
  wire  _GEN_21346 = _GEN_42097 | _GEN_19169; // @[rob.scala 145:{52,52}]
  wire  _GEN_21347 = _GEN_42098 | _GEN_19170; // @[rob.scala 145:{52,52}]
  wire  _GEN_21348 = _GEN_42099 | _GEN_19171; // @[rob.scala 145:{52,52}]
  wire  _GEN_21349 = _GEN_42100 | _GEN_19172; // @[rob.scala 145:{52,52}]
  wire  _GEN_21350 = _GEN_42101 | _GEN_19173; // @[rob.scala 145:{52,52}]
  wire  _GEN_21351 = _GEN_42102 | _GEN_19174; // @[rob.scala 145:{52,52}]
  wire  _GEN_21352 = _GEN_42103 | _GEN_19175; // @[rob.scala 145:{52,52}]
  wire  _GEN_21353 = _GEN_42104 | _GEN_19176; // @[rob.scala 145:{52,52}]
  wire  _GEN_21354 = _GEN_42105 | _GEN_19177; // @[rob.scala 145:{52,52}]
  wire  _GEN_21355 = _GEN_42106 | _GEN_19178; // @[rob.scala 145:{52,52}]
  wire  _GEN_21356 = _GEN_42107 | _GEN_19179; // @[rob.scala 145:{52,52}]
  wire  _GEN_21357 = _GEN_42108 | _GEN_19180; // @[rob.scala 145:{52,52}]
  wire  _GEN_21358 = _GEN_42109 | _GEN_19181; // @[rob.scala 145:{52,52}]
  wire  _GEN_21359 = _GEN_42110 | _GEN_19182; // @[rob.scala 145:{52,52}]
  wire  _GEN_21360 = _GEN_42111 | _GEN_19183; // @[rob.scala 145:{52,52}]
  wire  _GEN_21361 = _GEN_42112 | _GEN_19184; // @[rob.scala 145:{52,52}]
  wire  _GEN_21362 = _GEN_42113 | _GEN_19185; // @[rob.scala 145:{52,52}]
  wire  _GEN_21363 = _GEN_42114 | _GEN_19186; // @[rob.scala 145:{52,52}]
  wire  _GEN_21364 = _GEN_42115 | _GEN_19187; // @[rob.scala 145:{52,52}]
  wire  _GEN_21365 = _GEN_42116 | _GEN_19188; // @[rob.scala 145:{52,52}]
  wire  _GEN_21366 = _GEN_42117 | _GEN_19189; // @[rob.scala 145:{52,52}]
  wire  _GEN_21367 = _GEN_42118 | _GEN_19190; // @[rob.scala 145:{52,52}]
  wire  _GEN_21368 = _GEN_42119 | _GEN_19191; // @[rob.scala 145:{52,52}]
  wire  _GEN_21369 = _GEN_42120 | _GEN_19192; // @[rob.scala 145:{52,52}]
  wire  _GEN_21370 = _GEN_42121 | _GEN_19193; // @[rob.scala 145:{52,52}]
  wire  _GEN_21371 = _GEN_42122 | _GEN_19194; // @[rob.scala 145:{52,52}]
  wire  _GEN_21372 = _GEN_42123 | _GEN_19195; // @[rob.scala 145:{52,52}]
  wire  _GEN_21373 = _GEN_42124 | _GEN_19196; // @[rob.scala 145:{52,52}]
  wire  _GEN_21374 = _GEN_42125 | _GEN_19197; // @[rob.scala 145:{52,52}]
  wire  _GEN_21375 = _GEN_42126 | _GEN_19198; // @[rob.scala 145:{52,52}]
  wire  _GEN_21376 = _GEN_42127 | _GEN_19199; // @[rob.scala 145:{52,52}]
  wire  _GEN_21377 = _GEN_42128 | _GEN_19200; // @[rob.scala 145:{52,52}]
  wire  _GEN_21378 = io_i_ex_res_packs_0_valid ? _GEN_19202 : _GEN_19073; // @[rob.scala 141:39]
  wire  _GEN_21379 = io_i_ex_res_packs_0_valid ? _GEN_19203 : _GEN_19074; // @[rob.scala 141:39]
  wire  _GEN_21380 = io_i_ex_res_packs_0_valid ? _GEN_19204 : _GEN_19075; // @[rob.scala 141:39]
  wire  _GEN_21381 = io_i_ex_res_packs_0_valid ? _GEN_19205 : _GEN_19076; // @[rob.scala 141:39]
  wire  _GEN_21382 = io_i_ex_res_packs_0_valid ? _GEN_19206 : _GEN_19077; // @[rob.scala 141:39]
  wire  _GEN_21383 = io_i_ex_res_packs_0_valid ? _GEN_19207 : _GEN_19078; // @[rob.scala 141:39]
  wire  _GEN_21384 = io_i_ex_res_packs_0_valid ? _GEN_19208 : _GEN_19079; // @[rob.scala 141:39]
  wire  _GEN_21385 = io_i_ex_res_packs_0_valid ? _GEN_19209 : _GEN_19080; // @[rob.scala 141:39]
  wire  _GEN_21386 = io_i_ex_res_packs_0_valid ? _GEN_19210 : _GEN_19081; // @[rob.scala 141:39]
  wire  _GEN_21387 = io_i_ex_res_packs_0_valid ? _GEN_19211 : _GEN_19082; // @[rob.scala 141:39]
  wire  _GEN_21388 = io_i_ex_res_packs_0_valid ? _GEN_19212 : _GEN_19083; // @[rob.scala 141:39]
  wire  _GEN_21389 = io_i_ex_res_packs_0_valid ? _GEN_19213 : _GEN_19084; // @[rob.scala 141:39]
  wire  _GEN_21390 = io_i_ex_res_packs_0_valid ? _GEN_19214 : _GEN_19085; // @[rob.scala 141:39]
  wire  _GEN_21391 = io_i_ex_res_packs_0_valid ? _GEN_19215 : _GEN_19086; // @[rob.scala 141:39]
  wire  _GEN_21392 = io_i_ex_res_packs_0_valid ? _GEN_19216 : _GEN_19087; // @[rob.scala 141:39]
  wire  _GEN_21393 = io_i_ex_res_packs_0_valid ? _GEN_19217 : _GEN_19088; // @[rob.scala 141:39]
  wire  _GEN_21394 = io_i_ex_res_packs_0_valid ? _GEN_19218 : _GEN_19089; // @[rob.scala 141:39]
  wire  _GEN_21395 = io_i_ex_res_packs_0_valid ? _GEN_19219 : _GEN_19090; // @[rob.scala 141:39]
  wire  _GEN_21396 = io_i_ex_res_packs_0_valid ? _GEN_19220 : _GEN_19091; // @[rob.scala 141:39]
  wire  _GEN_21397 = io_i_ex_res_packs_0_valid ? _GEN_19221 : _GEN_19092; // @[rob.scala 141:39]
  wire  _GEN_21398 = io_i_ex_res_packs_0_valid ? _GEN_19222 : _GEN_19093; // @[rob.scala 141:39]
  wire  _GEN_21399 = io_i_ex_res_packs_0_valid ? _GEN_19223 : _GEN_19094; // @[rob.scala 141:39]
  wire  _GEN_21400 = io_i_ex_res_packs_0_valid ? _GEN_19224 : _GEN_19095; // @[rob.scala 141:39]
  wire  _GEN_21401 = io_i_ex_res_packs_0_valid ? _GEN_19225 : _GEN_19096; // @[rob.scala 141:39]
  wire  _GEN_21402 = io_i_ex_res_packs_0_valid ? _GEN_19226 : _GEN_19097; // @[rob.scala 141:39]
  wire  _GEN_21403 = io_i_ex_res_packs_0_valid ? _GEN_19227 : _GEN_19098; // @[rob.scala 141:39]
  wire  _GEN_21404 = io_i_ex_res_packs_0_valid ? _GEN_19228 : _GEN_19099; // @[rob.scala 141:39]
  wire  _GEN_21405 = io_i_ex_res_packs_0_valid ? _GEN_19229 : _GEN_19100; // @[rob.scala 141:39]
  wire  _GEN_21406 = io_i_ex_res_packs_0_valid ? _GEN_19230 : _GEN_19101; // @[rob.scala 141:39]
  wire  _GEN_21407 = io_i_ex_res_packs_0_valid ? _GEN_19231 : _GEN_19102; // @[rob.scala 141:39]
  wire  _GEN_21408 = io_i_ex_res_packs_0_valid ? _GEN_19232 : _GEN_19103; // @[rob.scala 141:39]
  wire  _GEN_21409 = io_i_ex_res_packs_0_valid ? _GEN_19233 : _GEN_19104; // @[rob.scala 141:39]
  wire  _GEN_21410 = io_i_ex_res_packs_0_valid ? _GEN_19234 : _GEN_19105; // @[rob.scala 141:39]
  wire  _GEN_21411 = io_i_ex_res_packs_0_valid ? _GEN_19235 : _GEN_19106; // @[rob.scala 141:39]
  wire  _GEN_21412 = io_i_ex_res_packs_0_valid ? _GEN_19236 : _GEN_19107; // @[rob.scala 141:39]
  wire  _GEN_21413 = io_i_ex_res_packs_0_valid ? _GEN_19237 : _GEN_19108; // @[rob.scala 141:39]
  wire  _GEN_21414 = io_i_ex_res_packs_0_valid ? _GEN_19238 : _GEN_19109; // @[rob.scala 141:39]
  wire  _GEN_21415 = io_i_ex_res_packs_0_valid ? _GEN_19239 : _GEN_19110; // @[rob.scala 141:39]
  wire  _GEN_21416 = io_i_ex_res_packs_0_valid ? _GEN_19240 : _GEN_19111; // @[rob.scala 141:39]
  wire  _GEN_21417 = io_i_ex_res_packs_0_valid ? _GEN_19241 : _GEN_19112; // @[rob.scala 141:39]
  wire  _GEN_21418 = io_i_ex_res_packs_0_valid ? _GEN_19242 : _GEN_19113; // @[rob.scala 141:39]
  wire  _GEN_21419 = io_i_ex_res_packs_0_valid ? _GEN_19243 : _GEN_19114; // @[rob.scala 141:39]
  wire  _GEN_21420 = io_i_ex_res_packs_0_valid ? _GEN_19244 : _GEN_19115; // @[rob.scala 141:39]
  wire  _GEN_21421 = io_i_ex_res_packs_0_valid ? _GEN_19245 : _GEN_19116; // @[rob.scala 141:39]
  wire  _GEN_21422 = io_i_ex_res_packs_0_valid ? _GEN_19246 : _GEN_19117; // @[rob.scala 141:39]
  wire  _GEN_21423 = io_i_ex_res_packs_0_valid ? _GEN_19247 : _GEN_19118; // @[rob.scala 141:39]
  wire  _GEN_21424 = io_i_ex_res_packs_0_valid ? _GEN_19248 : _GEN_19119; // @[rob.scala 141:39]
  wire  _GEN_21425 = io_i_ex_res_packs_0_valid ? _GEN_19249 : _GEN_19120; // @[rob.scala 141:39]
  wire  _GEN_21426 = io_i_ex_res_packs_0_valid ? _GEN_19250 : _GEN_19121; // @[rob.scala 141:39]
  wire  _GEN_21427 = io_i_ex_res_packs_0_valid ? _GEN_19251 : _GEN_19122; // @[rob.scala 141:39]
  wire  _GEN_21428 = io_i_ex_res_packs_0_valid ? _GEN_19252 : _GEN_19123; // @[rob.scala 141:39]
  wire  _GEN_21429 = io_i_ex_res_packs_0_valid ? _GEN_19253 : _GEN_19124; // @[rob.scala 141:39]
  wire  _GEN_21430 = io_i_ex_res_packs_0_valid ? _GEN_19254 : _GEN_19125; // @[rob.scala 141:39]
  wire  _GEN_21431 = io_i_ex_res_packs_0_valid ? _GEN_19255 : _GEN_19126; // @[rob.scala 141:39]
  wire  _GEN_21432 = io_i_ex_res_packs_0_valid ? _GEN_19256 : _GEN_19127; // @[rob.scala 141:39]
  wire  _GEN_21433 = io_i_ex_res_packs_0_valid ? _GEN_19257 : _GEN_19128; // @[rob.scala 141:39]
  wire  _GEN_21434 = io_i_ex_res_packs_0_valid ? _GEN_19258 : _GEN_19129; // @[rob.scala 141:39]
  wire  _GEN_21435 = io_i_ex_res_packs_0_valid ? _GEN_19259 : _GEN_19130; // @[rob.scala 141:39]
  wire  _GEN_21436 = io_i_ex_res_packs_0_valid ? _GEN_19260 : _GEN_19131; // @[rob.scala 141:39]
  wire  _GEN_21437 = io_i_ex_res_packs_0_valid ? _GEN_19261 : _GEN_19132; // @[rob.scala 141:39]
  wire  _GEN_21438 = io_i_ex_res_packs_0_valid ? _GEN_19262 : _GEN_19133; // @[rob.scala 141:39]
  wire  _GEN_21439 = io_i_ex_res_packs_0_valid ? _GEN_19263 : _GEN_19134; // @[rob.scala 141:39]
  wire  _GEN_21440 = io_i_ex_res_packs_0_valid ? _GEN_19264 : _GEN_19135; // @[rob.scala 141:39]
  wire  _GEN_21441 = io_i_ex_res_packs_0_valid ? _GEN_19265 : _GEN_19136; // @[rob.scala 141:39]
  wire [31:0] _GEN_21506 = io_i_ex_res_packs_0_valid ? _GEN_19330 : _GEN_17153; // @[rob.scala 141:39]
  wire [31:0] _GEN_21507 = io_i_ex_res_packs_0_valid ? _GEN_19331 : _GEN_17154; // @[rob.scala 141:39]
  wire [31:0] _GEN_21508 = io_i_ex_res_packs_0_valid ? _GEN_19332 : _GEN_17155; // @[rob.scala 141:39]
  wire [31:0] _GEN_21509 = io_i_ex_res_packs_0_valid ? _GEN_19333 : _GEN_17156; // @[rob.scala 141:39]
  wire [31:0] _GEN_21510 = io_i_ex_res_packs_0_valid ? _GEN_19334 : _GEN_17157; // @[rob.scala 141:39]
  wire [31:0] _GEN_21511 = io_i_ex_res_packs_0_valid ? _GEN_19335 : _GEN_17158; // @[rob.scala 141:39]
  wire [31:0] _GEN_21512 = io_i_ex_res_packs_0_valid ? _GEN_19336 : _GEN_17159; // @[rob.scala 141:39]
  wire [31:0] _GEN_21513 = io_i_ex_res_packs_0_valid ? _GEN_19337 : _GEN_17160; // @[rob.scala 141:39]
  wire [31:0] _GEN_21514 = io_i_ex_res_packs_0_valid ? _GEN_19338 : _GEN_17161; // @[rob.scala 141:39]
  wire [31:0] _GEN_21515 = io_i_ex_res_packs_0_valid ? _GEN_19339 : _GEN_17162; // @[rob.scala 141:39]
  wire [31:0] _GEN_21516 = io_i_ex_res_packs_0_valid ? _GEN_19340 : _GEN_17163; // @[rob.scala 141:39]
  wire [31:0] _GEN_21517 = io_i_ex_res_packs_0_valid ? _GEN_19341 : _GEN_17164; // @[rob.scala 141:39]
  wire [31:0] _GEN_21518 = io_i_ex_res_packs_0_valid ? _GEN_19342 : _GEN_17165; // @[rob.scala 141:39]
  wire [31:0] _GEN_21519 = io_i_ex_res_packs_0_valid ? _GEN_19343 : _GEN_17166; // @[rob.scala 141:39]
  wire [31:0] _GEN_21520 = io_i_ex_res_packs_0_valid ? _GEN_19344 : _GEN_17167; // @[rob.scala 141:39]
  wire [31:0] _GEN_21521 = io_i_ex_res_packs_0_valid ? _GEN_19345 : _GEN_17168; // @[rob.scala 141:39]
  wire [31:0] _GEN_21522 = io_i_ex_res_packs_0_valid ? _GEN_19346 : _GEN_17169; // @[rob.scala 141:39]
  wire [31:0] _GEN_21523 = io_i_ex_res_packs_0_valid ? _GEN_19347 : _GEN_17170; // @[rob.scala 141:39]
  wire [31:0] _GEN_21524 = io_i_ex_res_packs_0_valid ? _GEN_19348 : _GEN_17171; // @[rob.scala 141:39]
  wire [31:0] _GEN_21525 = io_i_ex_res_packs_0_valid ? _GEN_19349 : _GEN_17172; // @[rob.scala 141:39]
  wire [31:0] _GEN_21526 = io_i_ex_res_packs_0_valid ? _GEN_19350 : _GEN_17173; // @[rob.scala 141:39]
  wire [31:0] _GEN_21527 = io_i_ex_res_packs_0_valid ? _GEN_19351 : _GEN_17174; // @[rob.scala 141:39]
  wire [31:0] _GEN_21528 = io_i_ex_res_packs_0_valid ? _GEN_19352 : _GEN_17175; // @[rob.scala 141:39]
  wire [31:0] _GEN_21529 = io_i_ex_res_packs_0_valid ? _GEN_19353 : _GEN_17176; // @[rob.scala 141:39]
  wire [31:0] _GEN_21530 = io_i_ex_res_packs_0_valid ? _GEN_19354 : _GEN_17177; // @[rob.scala 141:39]
  wire [31:0] _GEN_21531 = io_i_ex_res_packs_0_valid ? _GEN_19355 : _GEN_17178; // @[rob.scala 141:39]
  wire [31:0] _GEN_21532 = io_i_ex_res_packs_0_valid ? _GEN_19356 : _GEN_17179; // @[rob.scala 141:39]
  wire [31:0] _GEN_21533 = io_i_ex_res_packs_0_valid ? _GEN_19357 : _GEN_17180; // @[rob.scala 141:39]
  wire [31:0] _GEN_21534 = io_i_ex_res_packs_0_valid ? _GEN_19358 : _GEN_17181; // @[rob.scala 141:39]
  wire [31:0] _GEN_21535 = io_i_ex_res_packs_0_valid ? _GEN_19359 : _GEN_17182; // @[rob.scala 141:39]
  wire [31:0] _GEN_21536 = io_i_ex_res_packs_0_valid ? _GEN_19360 : _GEN_17183; // @[rob.scala 141:39]
  wire [31:0] _GEN_21537 = io_i_ex_res_packs_0_valid ? _GEN_19361 : _GEN_17184; // @[rob.scala 141:39]
  wire [31:0] _GEN_21538 = io_i_ex_res_packs_0_valid ? _GEN_19362 : _GEN_17185; // @[rob.scala 141:39]
  wire [31:0] _GEN_21539 = io_i_ex_res_packs_0_valid ? _GEN_19363 : _GEN_17186; // @[rob.scala 141:39]
  wire [31:0] _GEN_21540 = io_i_ex_res_packs_0_valid ? _GEN_19364 : _GEN_17187; // @[rob.scala 141:39]
  wire [31:0] _GEN_21541 = io_i_ex_res_packs_0_valid ? _GEN_19365 : _GEN_17188; // @[rob.scala 141:39]
  wire [31:0] _GEN_21542 = io_i_ex_res_packs_0_valid ? _GEN_19366 : _GEN_17189; // @[rob.scala 141:39]
  wire [31:0] _GEN_21543 = io_i_ex_res_packs_0_valid ? _GEN_19367 : _GEN_17190; // @[rob.scala 141:39]
  wire [31:0] _GEN_21544 = io_i_ex_res_packs_0_valid ? _GEN_19368 : _GEN_17191; // @[rob.scala 141:39]
  wire [31:0] _GEN_21545 = io_i_ex_res_packs_0_valid ? _GEN_19369 : _GEN_17192; // @[rob.scala 141:39]
  wire [31:0] _GEN_21546 = io_i_ex_res_packs_0_valid ? _GEN_19370 : _GEN_17193; // @[rob.scala 141:39]
  wire [31:0] _GEN_21547 = io_i_ex_res_packs_0_valid ? _GEN_19371 : _GEN_17194; // @[rob.scala 141:39]
  wire [31:0] _GEN_21548 = io_i_ex_res_packs_0_valid ? _GEN_19372 : _GEN_17195; // @[rob.scala 141:39]
  wire [31:0] _GEN_21549 = io_i_ex_res_packs_0_valid ? _GEN_19373 : _GEN_17196; // @[rob.scala 141:39]
  wire [31:0] _GEN_21550 = io_i_ex_res_packs_0_valid ? _GEN_19374 : _GEN_17197; // @[rob.scala 141:39]
  wire [31:0] _GEN_21551 = io_i_ex_res_packs_0_valid ? _GEN_19375 : _GEN_17198; // @[rob.scala 141:39]
  wire [31:0] _GEN_21552 = io_i_ex_res_packs_0_valid ? _GEN_19376 : _GEN_17199; // @[rob.scala 141:39]
  wire [31:0] _GEN_21553 = io_i_ex_res_packs_0_valid ? _GEN_19377 : _GEN_17200; // @[rob.scala 141:39]
  wire [31:0] _GEN_21554 = io_i_ex_res_packs_0_valid ? _GEN_19378 : _GEN_17201; // @[rob.scala 141:39]
  wire [31:0] _GEN_21555 = io_i_ex_res_packs_0_valid ? _GEN_19379 : _GEN_17202; // @[rob.scala 141:39]
  wire [31:0] _GEN_21556 = io_i_ex_res_packs_0_valid ? _GEN_19380 : _GEN_17203; // @[rob.scala 141:39]
  wire [31:0] _GEN_21557 = io_i_ex_res_packs_0_valid ? _GEN_19381 : _GEN_17204; // @[rob.scala 141:39]
  wire [31:0] _GEN_21558 = io_i_ex_res_packs_0_valid ? _GEN_19382 : _GEN_17205; // @[rob.scala 141:39]
  wire [31:0] _GEN_21559 = io_i_ex_res_packs_0_valid ? _GEN_19383 : _GEN_17206; // @[rob.scala 141:39]
  wire [31:0] _GEN_21560 = io_i_ex_res_packs_0_valid ? _GEN_19384 : _GEN_17207; // @[rob.scala 141:39]
  wire [31:0] _GEN_21561 = io_i_ex_res_packs_0_valid ? _GEN_19385 : _GEN_17208; // @[rob.scala 141:39]
  wire [31:0] _GEN_21562 = io_i_ex_res_packs_0_valid ? _GEN_19386 : _GEN_17209; // @[rob.scala 141:39]
  wire [31:0] _GEN_21563 = io_i_ex_res_packs_0_valid ? _GEN_19387 : _GEN_17210; // @[rob.scala 141:39]
  wire [31:0] _GEN_21564 = io_i_ex_res_packs_0_valid ? _GEN_19388 : _GEN_17211; // @[rob.scala 141:39]
  wire [31:0] _GEN_21565 = io_i_ex_res_packs_0_valid ? _GEN_19389 : _GEN_17212; // @[rob.scala 141:39]
  wire [31:0] _GEN_21566 = io_i_ex_res_packs_0_valid ? _GEN_19390 : _GEN_17213; // @[rob.scala 141:39]
  wire [31:0] _GEN_21567 = io_i_ex_res_packs_0_valid ? _GEN_19391 : _GEN_17214; // @[rob.scala 141:39]
  wire [31:0] _GEN_21568 = io_i_ex_res_packs_0_valid ? _GEN_19392 : _GEN_17215; // @[rob.scala 141:39]
  wire [31:0] _GEN_21569 = io_i_ex_res_packs_0_valid ? _GEN_19393 : _GEN_17216; // @[rob.scala 141:39]
  wire [31:0] _GEN_21570 = io_i_ex_res_packs_0_valid ? _GEN_19394 : _GEN_17217; // @[rob.scala 141:39]
  wire [31:0] _GEN_21571 = io_i_ex_res_packs_0_valid ? _GEN_19395 : _GEN_17218; // @[rob.scala 141:39]
  wire [31:0] _GEN_21572 = io_i_ex_res_packs_0_valid ? _GEN_19396 : _GEN_17219; // @[rob.scala 141:39]
  wire [31:0] _GEN_21573 = io_i_ex_res_packs_0_valid ? _GEN_19397 : _GEN_17220; // @[rob.scala 141:39]
  wire [31:0] _GEN_21574 = io_i_ex_res_packs_0_valid ? _GEN_19398 : _GEN_17221; // @[rob.scala 141:39]
  wire [31:0] _GEN_21575 = io_i_ex_res_packs_0_valid ? _GEN_19399 : _GEN_17222; // @[rob.scala 141:39]
  wire [31:0] _GEN_21576 = io_i_ex_res_packs_0_valid ? _GEN_19400 : _GEN_17223; // @[rob.scala 141:39]
  wire [31:0] _GEN_21577 = io_i_ex_res_packs_0_valid ? _GEN_19401 : _GEN_17224; // @[rob.scala 141:39]
  wire [31:0] _GEN_21578 = io_i_ex_res_packs_0_valid ? _GEN_19402 : _GEN_17225; // @[rob.scala 141:39]
  wire [31:0] _GEN_21579 = io_i_ex_res_packs_0_valid ? _GEN_19403 : _GEN_17226; // @[rob.scala 141:39]
  wire [31:0] _GEN_21580 = io_i_ex_res_packs_0_valid ? _GEN_19404 : _GEN_17227; // @[rob.scala 141:39]
  wire [31:0] _GEN_21581 = io_i_ex_res_packs_0_valid ? _GEN_19405 : _GEN_17228; // @[rob.scala 141:39]
  wire [31:0] _GEN_21582 = io_i_ex_res_packs_0_valid ? _GEN_19406 : _GEN_17229; // @[rob.scala 141:39]
  wire [31:0] _GEN_21583 = io_i_ex_res_packs_0_valid ? _GEN_19407 : _GEN_17230; // @[rob.scala 141:39]
  wire [31:0] _GEN_21584 = io_i_ex_res_packs_0_valid ? _GEN_19408 : _GEN_17231; // @[rob.scala 141:39]
  wire [31:0] _GEN_21585 = io_i_ex_res_packs_0_valid ? _GEN_19409 : _GEN_17232; // @[rob.scala 141:39]
  wire [31:0] _GEN_21586 = io_i_ex_res_packs_0_valid ? _GEN_19410 : _GEN_17233; // @[rob.scala 141:39]
  wire [31:0] _GEN_21587 = io_i_ex_res_packs_0_valid ? _GEN_19411 : _GEN_17234; // @[rob.scala 141:39]
  wire [31:0] _GEN_21588 = io_i_ex_res_packs_0_valid ? _GEN_19412 : _GEN_17235; // @[rob.scala 141:39]
  wire [31:0] _GEN_21589 = io_i_ex_res_packs_0_valid ? _GEN_19413 : _GEN_17236; // @[rob.scala 141:39]
  wire [31:0] _GEN_21590 = io_i_ex_res_packs_0_valid ? _GEN_19414 : _GEN_17237; // @[rob.scala 141:39]
  wire [31:0] _GEN_21591 = io_i_ex_res_packs_0_valid ? _GEN_19415 : _GEN_17238; // @[rob.scala 141:39]
  wire [31:0] _GEN_21592 = io_i_ex_res_packs_0_valid ? _GEN_19416 : _GEN_17239; // @[rob.scala 141:39]
  wire [31:0] _GEN_21593 = io_i_ex_res_packs_0_valid ? _GEN_19417 : _GEN_17240; // @[rob.scala 141:39]
  wire [31:0] _GEN_21594 = io_i_ex_res_packs_0_valid ? _GEN_19418 : _GEN_17241; // @[rob.scala 141:39]
  wire [31:0] _GEN_21595 = io_i_ex_res_packs_0_valid ? _GEN_19419 : _GEN_17242; // @[rob.scala 141:39]
  wire [31:0] _GEN_21596 = io_i_ex_res_packs_0_valid ? _GEN_19420 : _GEN_17243; // @[rob.scala 141:39]
  wire [31:0] _GEN_21597 = io_i_ex_res_packs_0_valid ? _GEN_19421 : _GEN_17244; // @[rob.scala 141:39]
  wire [31:0] _GEN_21598 = io_i_ex_res_packs_0_valid ? _GEN_19422 : _GEN_17245; // @[rob.scala 141:39]
  wire [31:0] _GEN_21599 = io_i_ex_res_packs_0_valid ? _GEN_19423 : _GEN_17246; // @[rob.scala 141:39]
  wire [31:0] _GEN_21600 = io_i_ex_res_packs_0_valid ? _GEN_19424 : _GEN_17247; // @[rob.scala 141:39]
  wire [31:0] _GEN_21601 = io_i_ex_res_packs_0_valid ? _GEN_19425 : _GEN_17248; // @[rob.scala 141:39]
  wire [31:0] _GEN_21602 = io_i_ex_res_packs_0_valid ? _GEN_19426 : _GEN_17249; // @[rob.scala 141:39]
  wire [31:0] _GEN_21603 = io_i_ex_res_packs_0_valid ? _GEN_19427 : _GEN_17250; // @[rob.scala 141:39]
  wire [31:0] _GEN_21604 = io_i_ex_res_packs_0_valid ? _GEN_19428 : _GEN_17251; // @[rob.scala 141:39]
  wire [31:0] _GEN_21605 = io_i_ex_res_packs_0_valid ? _GEN_19429 : _GEN_17252; // @[rob.scala 141:39]
  wire [31:0] _GEN_21606 = io_i_ex_res_packs_0_valid ? _GEN_19430 : _GEN_17253; // @[rob.scala 141:39]
  wire [31:0] _GEN_21607 = io_i_ex_res_packs_0_valid ? _GEN_19431 : _GEN_17254; // @[rob.scala 141:39]
  wire [31:0] _GEN_21608 = io_i_ex_res_packs_0_valid ? _GEN_19432 : _GEN_17255; // @[rob.scala 141:39]
  wire [31:0] _GEN_21609 = io_i_ex_res_packs_0_valid ? _GEN_19433 : _GEN_17256; // @[rob.scala 141:39]
  wire [31:0] _GEN_21610 = io_i_ex_res_packs_0_valid ? _GEN_19434 : _GEN_17257; // @[rob.scala 141:39]
  wire [31:0] _GEN_21611 = io_i_ex_res_packs_0_valid ? _GEN_19435 : _GEN_17258; // @[rob.scala 141:39]
  wire [31:0] _GEN_21612 = io_i_ex_res_packs_0_valid ? _GEN_19436 : _GEN_17259; // @[rob.scala 141:39]
  wire [31:0] _GEN_21613 = io_i_ex_res_packs_0_valid ? _GEN_19437 : _GEN_17260; // @[rob.scala 141:39]
  wire [31:0] _GEN_21614 = io_i_ex_res_packs_0_valid ? _GEN_19438 : _GEN_17261; // @[rob.scala 141:39]
  wire [31:0] _GEN_21615 = io_i_ex_res_packs_0_valid ? _GEN_19439 : _GEN_17262; // @[rob.scala 141:39]
  wire [31:0] _GEN_21616 = io_i_ex_res_packs_0_valid ? _GEN_19440 : _GEN_17263; // @[rob.scala 141:39]
  wire [31:0] _GEN_21617 = io_i_ex_res_packs_0_valid ? _GEN_19441 : _GEN_17264; // @[rob.scala 141:39]
  wire [31:0] _GEN_21618 = io_i_ex_res_packs_0_valid ? _GEN_19442 : _GEN_17265; // @[rob.scala 141:39]
  wire [31:0] _GEN_21619 = io_i_ex_res_packs_0_valid ? _GEN_19443 : _GEN_17266; // @[rob.scala 141:39]
  wire [31:0] _GEN_21620 = io_i_ex_res_packs_0_valid ? _GEN_19444 : _GEN_17267; // @[rob.scala 141:39]
  wire [31:0] _GEN_21621 = io_i_ex_res_packs_0_valid ? _GEN_19445 : _GEN_17268; // @[rob.scala 141:39]
  wire [31:0] _GEN_21622 = io_i_ex_res_packs_0_valid ? _GEN_19446 : _GEN_17269; // @[rob.scala 141:39]
  wire [31:0] _GEN_21623 = io_i_ex_res_packs_0_valid ? _GEN_19447 : _GEN_17270; // @[rob.scala 141:39]
  wire [31:0] _GEN_21624 = io_i_ex_res_packs_0_valid ? _GEN_19448 : _GEN_17271; // @[rob.scala 141:39]
  wire [31:0] _GEN_21625 = io_i_ex_res_packs_0_valid ? _GEN_19449 : _GEN_17272; // @[rob.scala 141:39]
  wire [31:0] _GEN_21626 = io_i_ex_res_packs_0_valid ? _GEN_19450 : _GEN_17273; // @[rob.scala 141:39]
  wire [31:0] _GEN_21627 = io_i_ex_res_packs_0_valid ? _GEN_19451 : _GEN_17274; // @[rob.scala 141:39]
  wire [31:0] _GEN_21628 = io_i_ex_res_packs_0_valid ? _GEN_19452 : _GEN_17275; // @[rob.scala 141:39]
  wire [31:0] _GEN_21629 = io_i_ex_res_packs_0_valid ? _GEN_19453 : _GEN_17276; // @[rob.scala 141:39]
  wire [31:0] _GEN_21630 = io_i_ex_res_packs_0_valid ? _GEN_19454 : _GEN_17277; // @[rob.scala 141:39]
  wire [31:0] _GEN_21631 = io_i_ex_res_packs_0_valid ? _GEN_19455 : _GEN_17278; // @[rob.scala 141:39]
  wire [31:0] _GEN_21632 = io_i_ex_res_packs_0_valid ? _GEN_19456 : _GEN_17279; // @[rob.scala 141:39]
  wire [31:0] _GEN_21633 = io_i_ex_res_packs_0_valid ? _GEN_19457 : _GEN_17280; // @[rob.scala 141:39]
  wire [6:0] _GEN_21634 = io_i_ex_res_packs_0_valid ? _GEN_19458 : _GEN_17281; // @[rob.scala 141:39]
  wire [6:0] _GEN_21635 = io_i_ex_res_packs_0_valid ? _GEN_19459 : _GEN_17282; // @[rob.scala 141:39]
  wire [6:0] _GEN_21636 = io_i_ex_res_packs_0_valid ? _GEN_19460 : _GEN_17283; // @[rob.scala 141:39]
  wire [6:0] _GEN_21637 = io_i_ex_res_packs_0_valid ? _GEN_19461 : _GEN_17284; // @[rob.scala 141:39]
  wire [6:0] _GEN_21638 = io_i_ex_res_packs_0_valid ? _GEN_19462 : _GEN_17285; // @[rob.scala 141:39]
  wire [6:0] _GEN_21639 = io_i_ex_res_packs_0_valid ? _GEN_19463 : _GEN_17286; // @[rob.scala 141:39]
  wire [6:0] _GEN_21640 = io_i_ex_res_packs_0_valid ? _GEN_19464 : _GEN_17287; // @[rob.scala 141:39]
  wire [6:0] _GEN_21641 = io_i_ex_res_packs_0_valid ? _GEN_19465 : _GEN_17288; // @[rob.scala 141:39]
  wire [6:0] _GEN_21642 = io_i_ex_res_packs_0_valid ? _GEN_19466 : _GEN_17289; // @[rob.scala 141:39]
  wire [6:0] _GEN_21643 = io_i_ex_res_packs_0_valid ? _GEN_19467 : _GEN_17290; // @[rob.scala 141:39]
  wire [6:0] _GEN_21644 = io_i_ex_res_packs_0_valid ? _GEN_19468 : _GEN_17291; // @[rob.scala 141:39]
  wire [6:0] _GEN_21645 = io_i_ex_res_packs_0_valid ? _GEN_19469 : _GEN_17292; // @[rob.scala 141:39]
  wire [6:0] _GEN_21646 = io_i_ex_res_packs_0_valid ? _GEN_19470 : _GEN_17293; // @[rob.scala 141:39]
  wire [6:0] _GEN_21647 = io_i_ex_res_packs_0_valid ? _GEN_19471 : _GEN_17294; // @[rob.scala 141:39]
  wire [6:0] _GEN_21648 = io_i_ex_res_packs_0_valid ? _GEN_19472 : _GEN_17295; // @[rob.scala 141:39]
  wire [6:0] _GEN_21649 = io_i_ex_res_packs_0_valid ? _GEN_19473 : _GEN_17296; // @[rob.scala 141:39]
  wire [6:0] _GEN_21650 = io_i_ex_res_packs_0_valid ? _GEN_19474 : _GEN_17297; // @[rob.scala 141:39]
  wire [6:0] _GEN_21651 = io_i_ex_res_packs_0_valid ? _GEN_19475 : _GEN_17298; // @[rob.scala 141:39]
  wire [6:0] _GEN_21652 = io_i_ex_res_packs_0_valid ? _GEN_19476 : _GEN_17299; // @[rob.scala 141:39]
  wire [6:0] _GEN_21653 = io_i_ex_res_packs_0_valid ? _GEN_19477 : _GEN_17300; // @[rob.scala 141:39]
  wire [6:0] _GEN_21654 = io_i_ex_res_packs_0_valid ? _GEN_19478 : _GEN_17301; // @[rob.scala 141:39]
  wire [6:0] _GEN_21655 = io_i_ex_res_packs_0_valid ? _GEN_19479 : _GEN_17302; // @[rob.scala 141:39]
  wire [6:0] _GEN_21656 = io_i_ex_res_packs_0_valid ? _GEN_19480 : _GEN_17303; // @[rob.scala 141:39]
  wire [6:0] _GEN_21657 = io_i_ex_res_packs_0_valid ? _GEN_19481 : _GEN_17304; // @[rob.scala 141:39]
  wire [6:0] _GEN_21658 = io_i_ex_res_packs_0_valid ? _GEN_19482 : _GEN_17305; // @[rob.scala 141:39]
  wire [6:0] _GEN_21659 = io_i_ex_res_packs_0_valid ? _GEN_19483 : _GEN_17306; // @[rob.scala 141:39]
  wire [6:0] _GEN_21660 = io_i_ex_res_packs_0_valid ? _GEN_19484 : _GEN_17307; // @[rob.scala 141:39]
  wire [6:0] _GEN_21661 = io_i_ex_res_packs_0_valid ? _GEN_19485 : _GEN_17308; // @[rob.scala 141:39]
  wire [6:0] _GEN_21662 = io_i_ex_res_packs_0_valid ? _GEN_19486 : _GEN_17309; // @[rob.scala 141:39]
  wire [6:0] _GEN_21663 = io_i_ex_res_packs_0_valid ? _GEN_19487 : _GEN_17310; // @[rob.scala 141:39]
  wire [6:0] _GEN_21664 = io_i_ex_res_packs_0_valid ? _GEN_19488 : _GEN_17311; // @[rob.scala 141:39]
  wire [6:0] _GEN_21665 = io_i_ex_res_packs_0_valid ? _GEN_19489 : _GEN_17312; // @[rob.scala 141:39]
  wire [6:0] _GEN_21666 = io_i_ex_res_packs_0_valid ? _GEN_19490 : _GEN_17313; // @[rob.scala 141:39]
  wire [6:0] _GEN_21667 = io_i_ex_res_packs_0_valid ? _GEN_19491 : _GEN_17314; // @[rob.scala 141:39]
  wire [6:0] _GEN_21668 = io_i_ex_res_packs_0_valid ? _GEN_19492 : _GEN_17315; // @[rob.scala 141:39]
  wire [6:0] _GEN_21669 = io_i_ex_res_packs_0_valid ? _GEN_19493 : _GEN_17316; // @[rob.scala 141:39]
  wire [6:0] _GEN_21670 = io_i_ex_res_packs_0_valid ? _GEN_19494 : _GEN_17317; // @[rob.scala 141:39]
  wire [6:0] _GEN_21671 = io_i_ex_res_packs_0_valid ? _GEN_19495 : _GEN_17318; // @[rob.scala 141:39]
  wire [6:0] _GEN_21672 = io_i_ex_res_packs_0_valid ? _GEN_19496 : _GEN_17319; // @[rob.scala 141:39]
  wire [6:0] _GEN_21673 = io_i_ex_res_packs_0_valid ? _GEN_19497 : _GEN_17320; // @[rob.scala 141:39]
  wire [6:0] _GEN_21674 = io_i_ex_res_packs_0_valid ? _GEN_19498 : _GEN_17321; // @[rob.scala 141:39]
  wire [6:0] _GEN_21675 = io_i_ex_res_packs_0_valid ? _GEN_19499 : _GEN_17322; // @[rob.scala 141:39]
  wire [6:0] _GEN_21676 = io_i_ex_res_packs_0_valid ? _GEN_19500 : _GEN_17323; // @[rob.scala 141:39]
  wire [6:0] _GEN_21677 = io_i_ex_res_packs_0_valid ? _GEN_19501 : _GEN_17324; // @[rob.scala 141:39]
  wire [6:0] _GEN_21678 = io_i_ex_res_packs_0_valid ? _GEN_19502 : _GEN_17325; // @[rob.scala 141:39]
  wire [6:0] _GEN_21679 = io_i_ex_res_packs_0_valid ? _GEN_19503 : _GEN_17326; // @[rob.scala 141:39]
  wire [6:0] _GEN_21680 = io_i_ex_res_packs_0_valid ? _GEN_19504 : _GEN_17327; // @[rob.scala 141:39]
  wire [6:0] _GEN_21681 = io_i_ex_res_packs_0_valid ? _GEN_19505 : _GEN_17328; // @[rob.scala 141:39]
  wire [6:0] _GEN_21682 = io_i_ex_res_packs_0_valid ? _GEN_19506 : _GEN_17329; // @[rob.scala 141:39]
  wire [6:0] _GEN_21683 = io_i_ex_res_packs_0_valid ? _GEN_19507 : _GEN_17330; // @[rob.scala 141:39]
  wire [6:0] _GEN_21684 = io_i_ex_res_packs_0_valid ? _GEN_19508 : _GEN_17331; // @[rob.scala 141:39]
  wire [6:0] _GEN_21685 = io_i_ex_res_packs_0_valid ? _GEN_19509 : _GEN_17332; // @[rob.scala 141:39]
  wire [6:0] _GEN_21686 = io_i_ex_res_packs_0_valid ? _GEN_19510 : _GEN_17333; // @[rob.scala 141:39]
  wire [6:0] _GEN_21687 = io_i_ex_res_packs_0_valid ? _GEN_19511 : _GEN_17334; // @[rob.scala 141:39]
  wire [6:0] _GEN_21688 = io_i_ex_res_packs_0_valid ? _GEN_19512 : _GEN_17335; // @[rob.scala 141:39]
  wire [6:0] _GEN_21689 = io_i_ex_res_packs_0_valid ? _GEN_19513 : _GEN_17336; // @[rob.scala 141:39]
  wire [6:0] _GEN_21690 = io_i_ex_res_packs_0_valid ? _GEN_19514 : _GEN_17337; // @[rob.scala 141:39]
  wire [6:0] _GEN_21691 = io_i_ex_res_packs_0_valid ? _GEN_19515 : _GEN_17338; // @[rob.scala 141:39]
  wire [6:0] _GEN_21692 = io_i_ex_res_packs_0_valid ? _GEN_19516 : _GEN_17339; // @[rob.scala 141:39]
  wire [6:0] _GEN_21693 = io_i_ex_res_packs_0_valid ? _GEN_19517 : _GEN_17340; // @[rob.scala 141:39]
  wire [6:0] _GEN_21694 = io_i_ex_res_packs_0_valid ? _GEN_19518 : _GEN_17341; // @[rob.scala 141:39]
  wire [6:0] _GEN_21695 = io_i_ex_res_packs_0_valid ? _GEN_19519 : _GEN_17342; // @[rob.scala 141:39]
  wire [6:0] _GEN_21696 = io_i_ex_res_packs_0_valid ? _GEN_19520 : _GEN_17343; // @[rob.scala 141:39]
  wire [6:0] _GEN_21697 = io_i_ex_res_packs_0_valid ? _GEN_19521 : _GEN_17344; // @[rob.scala 141:39]
  wire [6:0] _GEN_22018 = io_i_ex_res_packs_0_valid ? _GEN_19842 : _GEN_17665; // @[rob.scala 141:39]
  wire [6:0] _GEN_22019 = io_i_ex_res_packs_0_valid ? _GEN_19843 : _GEN_17666; // @[rob.scala 141:39]
  wire [6:0] _GEN_22020 = io_i_ex_res_packs_0_valid ? _GEN_19844 : _GEN_17667; // @[rob.scala 141:39]
  wire [6:0] _GEN_22021 = io_i_ex_res_packs_0_valid ? _GEN_19845 : _GEN_17668; // @[rob.scala 141:39]
  wire [6:0] _GEN_22022 = io_i_ex_res_packs_0_valid ? _GEN_19846 : _GEN_17669; // @[rob.scala 141:39]
  wire [6:0] _GEN_22023 = io_i_ex_res_packs_0_valid ? _GEN_19847 : _GEN_17670; // @[rob.scala 141:39]
  wire [6:0] _GEN_22024 = io_i_ex_res_packs_0_valid ? _GEN_19848 : _GEN_17671; // @[rob.scala 141:39]
  wire [6:0] _GEN_22025 = io_i_ex_res_packs_0_valid ? _GEN_19849 : _GEN_17672; // @[rob.scala 141:39]
  wire [6:0] _GEN_22026 = io_i_ex_res_packs_0_valid ? _GEN_19850 : _GEN_17673; // @[rob.scala 141:39]
  wire [6:0] _GEN_22027 = io_i_ex_res_packs_0_valid ? _GEN_19851 : _GEN_17674; // @[rob.scala 141:39]
  wire [6:0] _GEN_22028 = io_i_ex_res_packs_0_valid ? _GEN_19852 : _GEN_17675; // @[rob.scala 141:39]
  wire [6:0] _GEN_22029 = io_i_ex_res_packs_0_valid ? _GEN_19853 : _GEN_17676; // @[rob.scala 141:39]
  wire [6:0] _GEN_22030 = io_i_ex_res_packs_0_valid ? _GEN_19854 : _GEN_17677; // @[rob.scala 141:39]
  wire [6:0] _GEN_22031 = io_i_ex_res_packs_0_valid ? _GEN_19855 : _GEN_17678; // @[rob.scala 141:39]
  wire [6:0] _GEN_22032 = io_i_ex_res_packs_0_valid ? _GEN_19856 : _GEN_17679; // @[rob.scala 141:39]
  wire [6:0] _GEN_22033 = io_i_ex_res_packs_0_valid ? _GEN_19857 : _GEN_17680; // @[rob.scala 141:39]
  wire [6:0] _GEN_22034 = io_i_ex_res_packs_0_valid ? _GEN_19858 : _GEN_17681; // @[rob.scala 141:39]
  wire [6:0] _GEN_22035 = io_i_ex_res_packs_0_valid ? _GEN_19859 : _GEN_17682; // @[rob.scala 141:39]
  wire [6:0] _GEN_22036 = io_i_ex_res_packs_0_valid ? _GEN_19860 : _GEN_17683; // @[rob.scala 141:39]
  wire [6:0] _GEN_22037 = io_i_ex_res_packs_0_valid ? _GEN_19861 : _GEN_17684; // @[rob.scala 141:39]
  wire [6:0] _GEN_22038 = io_i_ex_res_packs_0_valid ? _GEN_19862 : _GEN_17685; // @[rob.scala 141:39]
  wire [6:0] _GEN_22039 = io_i_ex_res_packs_0_valid ? _GEN_19863 : _GEN_17686; // @[rob.scala 141:39]
  wire [6:0] _GEN_22040 = io_i_ex_res_packs_0_valid ? _GEN_19864 : _GEN_17687; // @[rob.scala 141:39]
  wire [6:0] _GEN_22041 = io_i_ex_res_packs_0_valid ? _GEN_19865 : _GEN_17688; // @[rob.scala 141:39]
  wire [6:0] _GEN_22042 = io_i_ex_res_packs_0_valid ? _GEN_19866 : _GEN_17689; // @[rob.scala 141:39]
  wire [6:0] _GEN_22043 = io_i_ex_res_packs_0_valid ? _GEN_19867 : _GEN_17690; // @[rob.scala 141:39]
  wire [6:0] _GEN_22044 = io_i_ex_res_packs_0_valid ? _GEN_19868 : _GEN_17691; // @[rob.scala 141:39]
  wire [6:0] _GEN_22045 = io_i_ex_res_packs_0_valid ? _GEN_19869 : _GEN_17692; // @[rob.scala 141:39]
  wire [6:0] _GEN_22046 = io_i_ex_res_packs_0_valid ? _GEN_19870 : _GEN_17693; // @[rob.scala 141:39]
  wire [6:0] _GEN_22047 = io_i_ex_res_packs_0_valid ? _GEN_19871 : _GEN_17694; // @[rob.scala 141:39]
  wire [6:0] _GEN_22048 = io_i_ex_res_packs_0_valid ? _GEN_19872 : _GEN_17695; // @[rob.scala 141:39]
  wire [6:0] _GEN_22049 = io_i_ex_res_packs_0_valid ? _GEN_19873 : _GEN_17696; // @[rob.scala 141:39]
  wire [6:0] _GEN_22050 = io_i_ex_res_packs_0_valid ? _GEN_19874 : _GEN_17697; // @[rob.scala 141:39]
  wire [6:0] _GEN_22051 = io_i_ex_res_packs_0_valid ? _GEN_19875 : _GEN_17698; // @[rob.scala 141:39]
  wire [6:0] _GEN_22052 = io_i_ex_res_packs_0_valid ? _GEN_19876 : _GEN_17699; // @[rob.scala 141:39]
  wire [6:0] _GEN_22053 = io_i_ex_res_packs_0_valid ? _GEN_19877 : _GEN_17700; // @[rob.scala 141:39]
  wire [6:0] _GEN_22054 = io_i_ex_res_packs_0_valid ? _GEN_19878 : _GEN_17701; // @[rob.scala 141:39]
  wire [6:0] _GEN_22055 = io_i_ex_res_packs_0_valid ? _GEN_19879 : _GEN_17702; // @[rob.scala 141:39]
  wire [6:0] _GEN_22056 = io_i_ex_res_packs_0_valid ? _GEN_19880 : _GEN_17703; // @[rob.scala 141:39]
  wire [6:0] _GEN_22057 = io_i_ex_res_packs_0_valid ? _GEN_19881 : _GEN_17704; // @[rob.scala 141:39]
  wire [6:0] _GEN_22058 = io_i_ex_res_packs_0_valid ? _GEN_19882 : _GEN_17705; // @[rob.scala 141:39]
  wire [6:0] _GEN_22059 = io_i_ex_res_packs_0_valid ? _GEN_19883 : _GEN_17706; // @[rob.scala 141:39]
  wire [6:0] _GEN_22060 = io_i_ex_res_packs_0_valid ? _GEN_19884 : _GEN_17707; // @[rob.scala 141:39]
  wire [6:0] _GEN_22061 = io_i_ex_res_packs_0_valid ? _GEN_19885 : _GEN_17708; // @[rob.scala 141:39]
  wire [6:0] _GEN_22062 = io_i_ex_res_packs_0_valid ? _GEN_19886 : _GEN_17709; // @[rob.scala 141:39]
  wire [6:0] _GEN_22063 = io_i_ex_res_packs_0_valid ? _GEN_19887 : _GEN_17710; // @[rob.scala 141:39]
  wire [6:0] _GEN_22064 = io_i_ex_res_packs_0_valid ? _GEN_19888 : _GEN_17711; // @[rob.scala 141:39]
  wire [6:0] _GEN_22065 = io_i_ex_res_packs_0_valid ? _GEN_19889 : _GEN_17712; // @[rob.scala 141:39]
  wire [6:0] _GEN_22066 = io_i_ex_res_packs_0_valid ? _GEN_19890 : _GEN_17713; // @[rob.scala 141:39]
  wire [6:0] _GEN_22067 = io_i_ex_res_packs_0_valid ? _GEN_19891 : _GEN_17714; // @[rob.scala 141:39]
  wire [6:0] _GEN_22068 = io_i_ex_res_packs_0_valid ? _GEN_19892 : _GEN_17715; // @[rob.scala 141:39]
  wire [6:0] _GEN_22069 = io_i_ex_res_packs_0_valid ? _GEN_19893 : _GEN_17716; // @[rob.scala 141:39]
  wire [6:0] _GEN_22070 = io_i_ex_res_packs_0_valid ? _GEN_19894 : _GEN_17717; // @[rob.scala 141:39]
  wire [6:0] _GEN_22071 = io_i_ex_res_packs_0_valid ? _GEN_19895 : _GEN_17718; // @[rob.scala 141:39]
  wire [6:0] _GEN_22072 = io_i_ex_res_packs_0_valid ? _GEN_19896 : _GEN_17719; // @[rob.scala 141:39]
  wire [6:0] _GEN_22073 = io_i_ex_res_packs_0_valid ? _GEN_19897 : _GEN_17720; // @[rob.scala 141:39]
  wire [6:0] _GEN_22074 = io_i_ex_res_packs_0_valid ? _GEN_19898 : _GEN_17721; // @[rob.scala 141:39]
  wire [6:0] _GEN_22075 = io_i_ex_res_packs_0_valid ? _GEN_19899 : _GEN_17722; // @[rob.scala 141:39]
  wire [6:0] _GEN_22076 = io_i_ex_res_packs_0_valid ? _GEN_19900 : _GEN_17723; // @[rob.scala 141:39]
  wire [6:0] _GEN_22077 = io_i_ex_res_packs_0_valid ? _GEN_19901 : _GEN_17724; // @[rob.scala 141:39]
  wire [6:0] _GEN_22078 = io_i_ex_res_packs_0_valid ? _GEN_19902 : _GEN_17725; // @[rob.scala 141:39]
  wire [6:0] _GEN_22079 = io_i_ex_res_packs_0_valid ? _GEN_19903 : _GEN_17726; // @[rob.scala 141:39]
  wire [6:0] _GEN_22080 = io_i_ex_res_packs_0_valid ? _GEN_19904 : _GEN_17727; // @[rob.scala 141:39]
  wire [6:0] _GEN_22081 = io_i_ex_res_packs_0_valid ? _GEN_19905 : _GEN_17728; // @[rob.scala 141:39]
  wire [6:0] _GEN_22082 = io_i_ex_res_packs_0_valid ? _GEN_19906 : _GEN_17729; // @[rob.scala 141:39]
  wire [6:0] _GEN_22083 = io_i_ex_res_packs_0_valid ? _GEN_19907 : _GEN_17730; // @[rob.scala 141:39]
  wire [6:0] _GEN_22084 = io_i_ex_res_packs_0_valid ? _GEN_19908 : _GEN_17731; // @[rob.scala 141:39]
  wire [6:0] _GEN_22085 = io_i_ex_res_packs_0_valid ? _GEN_19909 : _GEN_17732; // @[rob.scala 141:39]
  wire [6:0] _GEN_22086 = io_i_ex_res_packs_0_valid ? _GEN_19910 : _GEN_17733; // @[rob.scala 141:39]
  wire [6:0] _GEN_22087 = io_i_ex_res_packs_0_valid ? _GEN_19911 : _GEN_17734; // @[rob.scala 141:39]
  wire [6:0] _GEN_22088 = io_i_ex_res_packs_0_valid ? _GEN_19912 : _GEN_17735; // @[rob.scala 141:39]
  wire [6:0] _GEN_22089 = io_i_ex_res_packs_0_valid ? _GEN_19913 : _GEN_17736; // @[rob.scala 141:39]
  wire [6:0] _GEN_22090 = io_i_ex_res_packs_0_valid ? _GEN_19914 : _GEN_17737; // @[rob.scala 141:39]
  wire [6:0] _GEN_22091 = io_i_ex_res_packs_0_valid ? _GEN_19915 : _GEN_17738; // @[rob.scala 141:39]
  wire [6:0] _GEN_22092 = io_i_ex_res_packs_0_valid ? _GEN_19916 : _GEN_17739; // @[rob.scala 141:39]
  wire [6:0] _GEN_22093 = io_i_ex_res_packs_0_valid ? _GEN_19917 : _GEN_17740; // @[rob.scala 141:39]
  wire [6:0] _GEN_22094 = io_i_ex_res_packs_0_valid ? _GEN_19918 : _GEN_17741; // @[rob.scala 141:39]
  wire [6:0] _GEN_22095 = io_i_ex_res_packs_0_valid ? _GEN_19919 : _GEN_17742; // @[rob.scala 141:39]
  wire [6:0] _GEN_22096 = io_i_ex_res_packs_0_valid ? _GEN_19920 : _GEN_17743; // @[rob.scala 141:39]
  wire [6:0] _GEN_22097 = io_i_ex_res_packs_0_valid ? _GEN_19921 : _GEN_17744; // @[rob.scala 141:39]
  wire [6:0] _GEN_22098 = io_i_ex_res_packs_0_valid ? _GEN_19922 : _GEN_17745; // @[rob.scala 141:39]
  wire [6:0] _GEN_22099 = io_i_ex_res_packs_0_valid ? _GEN_19923 : _GEN_17746; // @[rob.scala 141:39]
  wire [6:0] _GEN_22100 = io_i_ex_res_packs_0_valid ? _GEN_19924 : _GEN_17747; // @[rob.scala 141:39]
  wire [6:0] _GEN_22101 = io_i_ex_res_packs_0_valid ? _GEN_19925 : _GEN_17748; // @[rob.scala 141:39]
  wire [6:0] _GEN_22102 = io_i_ex_res_packs_0_valid ? _GEN_19926 : _GEN_17749; // @[rob.scala 141:39]
  wire [6:0] _GEN_22103 = io_i_ex_res_packs_0_valid ? _GEN_19927 : _GEN_17750; // @[rob.scala 141:39]
  wire [6:0] _GEN_22104 = io_i_ex_res_packs_0_valid ? _GEN_19928 : _GEN_17751; // @[rob.scala 141:39]
  wire [6:0] _GEN_22105 = io_i_ex_res_packs_0_valid ? _GEN_19929 : _GEN_17752; // @[rob.scala 141:39]
  wire [6:0] _GEN_22106 = io_i_ex_res_packs_0_valid ? _GEN_19930 : _GEN_17753; // @[rob.scala 141:39]
  wire [6:0] _GEN_22107 = io_i_ex_res_packs_0_valid ? _GEN_19931 : _GEN_17754; // @[rob.scala 141:39]
  wire [6:0] _GEN_22108 = io_i_ex_res_packs_0_valid ? _GEN_19932 : _GEN_17755; // @[rob.scala 141:39]
  wire [6:0] _GEN_22109 = io_i_ex_res_packs_0_valid ? _GEN_19933 : _GEN_17756; // @[rob.scala 141:39]
  wire [6:0] _GEN_22110 = io_i_ex_res_packs_0_valid ? _GEN_19934 : _GEN_17757; // @[rob.scala 141:39]
  wire [6:0] _GEN_22111 = io_i_ex_res_packs_0_valid ? _GEN_19935 : _GEN_17758; // @[rob.scala 141:39]
  wire [6:0] _GEN_22112 = io_i_ex_res_packs_0_valid ? _GEN_19936 : _GEN_17759; // @[rob.scala 141:39]
  wire [6:0] _GEN_22113 = io_i_ex_res_packs_0_valid ? _GEN_19937 : _GEN_17760; // @[rob.scala 141:39]
  wire [6:0] _GEN_22114 = io_i_ex_res_packs_0_valid ? _GEN_19938 : _GEN_17761; // @[rob.scala 141:39]
  wire [6:0] _GEN_22115 = io_i_ex_res_packs_0_valid ? _GEN_19939 : _GEN_17762; // @[rob.scala 141:39]
  wire [6:0] _GEN_22116 = io_i_ex_res_packs_0_valid ? _GEN_19940 : _GEN_17763; // @[rob.scala 141:39]
  wire [6:0] _GEN_22117 = io_i_ex_res_packs_0_valid ? _GEN_19941 : _GEN_17764; // @[rob.scala 141:39]
  wire [6:0] _GEN_22118 = io_i_ex_res_packs_0_valid ? _GEN_19942 : _GEN_17765; // @[rob.scala 141:39]
  wire [6:0] _GEN_22119 = io_i_ex_res_packs_0_valid ? _GEN_19943 : _GEN_17766; // @[rob.scala 141:39]
  wire [6:0] _GEN_22120 = io_i_ex_res_packs_0_valid ? _GEN_19944 : _GEN_17767; // @[rob.scala 141:39]
  wire [6:0] _GEN_22121 = io_i_ex_res_packs_0_valid ? _GEN_19945 : _GEN_17768; // @[rob.scala 141:39]
  wire [6:0] _GEN_22122 = io_i_ex_res_packs_0_valid ? _GEN_19946 : _GEN_17769; // @[rob.scala 141:39]
  wire [6:0] _GEN_22123 = io_i_ex_res_packs_0_valid ? _GEN_19947 : _GEN_17770; // @[rob.scala 141:39]
  wire [6:0] _GEN_22124 = io_i_ex_res_packs_0_valid ? _GEN_19948 : _GEN_17771; // @[rob.scala 141:39]
  wire [6:0] _GEN_22125 = io_i_ex_res_packs_0_valid ? _GEN_19949 : _GEN_17772; // @[rob.scala 141:39]
  wire [6:0] _GEN_22126 = io_i_ex_res_packs_0_valid ? _GEN_19950 : _GEN_17773; // @[rob.scala 141:39]
  wire [6:0] _GEN_22127 = io_i_ex_res_packs_0_valid ? _GEN_19951 : _GEN_17774; // @[rob.scala 141:39]
  wire [6:0] _GEN_22128 = io_i_ex_res_packs_0_valid ? _GEN_19952 : _GEN_17775; // @[rob.scala 141:39]
  wire [6:0] _GEN_22129 = io_i_ex_res_packs_0_valid ? _GEN_19953 : _GEN_17776; // @[rob.scala 141:39]
  wire [6:0] _GEN_22130 = io_i_ex_res_packs_0_valid ? _GEN_19954 : _GEN_17777; // @[rob.scala 141:39]
  wire [6:0] _GEN_22131 = io_i_ex_res_packs_0_valid ? _GEN_19955 : _GEN_17778; // @[rob.scala 141:39]
  wire [6:0] _GEN_22132 = io_i_ex_res_packs_0_valid ? _GEN_19956 : _GEN_17779; // @[rob.scala 141:39]
  wire [6:0] _GEN_22133 = io_i_ex_res_packs_0_valid ? _GEN_19957 : _GEN_17780; // @[rob.scala 141:39]
  wire [6:0] _GEN_22134 = io_i_ex_res_packs_0_valid ? _GEN_19958 : _GEN_17781; // @[rob.scala 141:39]
  wire [6:0] _GEN_22135 = io_i_ex_res_packs_0_valid ? _GEN_19959 : _GEN_17782; // @[rob.scala 141:39]
  wire [6:0] _GEN_22136 = io_i_ex_res_packs_0_valid ? _GEN_19960 : _GEN_17783; // @[rob.scala 141:39]
  wire [6:0] _GEN_22137 = io_i_ex_res_packs_0_valid ? _GEN_19961 : _GEN_17784; // @[rob.scala 141:39]
  wire [6:0] _GEN_22138 = io_i_ex_res_packs_0_valid ? _GEN_19962 : _GEN_17785; // @[rob.scala 141:39]
  wire [6:0] _GEN_22139 = io_i_ex_res_packs_0_valid ? _GEN_19963 : _GEN_17786; // @[rob.scala 141:39]
  wire [6:0] _GEN_22140 = io_i_ex_res_packs_0_valid ? _GEN_19964 : _GEN_17787; // @[rob.scala 141:39]
  wire [6:0] _GEN_22141 = io_i_ex_res_packs_0_valid ? _GEN_19965 : _GEN_17788; // @[rob.scala 141:39]
  wire [6:0] _GEN_22142 = io_i_ex_res_packs_0_valid ? _GEN_19966 : _GEN_17789; // @[rob.scala 141:39]
  wire [6:0] _GEN_22143 = io_i_ex_res_packs_0_valid ? _GEN_19967 : _GEN_17790; // @[rob.scala 141:39]
  wire [6:0] _GEN_22144 = io_i_ex_res_packs_0_valid ? _GEN_19968 : _GEN_17791; // @[rob.scala 141:39]
  wire [6:0] _GEN_22145 = io_i_ex_res_packs_0_valid ? _GEN_19969 : _GEN_17792; // @[rob.scala 141:39]
  wire [4:0] _GEN_22146 = io_i_ex_res_packs_0_valid ? _GEN_19970 : _GEN_17793; // @[rob.scala 141:39]
  wire [4:0] _GEN_22147 = io_i_ex_res_packs_0_valid ? _GEN_19971 : _GEN_17794; // @[rob.scala 141:39]
  wire [4:0] _GEN_22148 = io_i_ex_res_packs_0_valid ? _GEN_19972 : _GEN_17795; // @[rob.scala 141:39]
  wire [4:0] _GEN_22149 = io_i_ex_res_packs_0_valid ? _GEN_19973 : _GEN_17796; // @[rob.scala 141:39]
  wire [4:0] _GEN_22150 = io_i_ex_res_packs_0_valid ? _GEN_19974 : _GEN_17797; // @[rob.scala 141:39]
  wire [4:0] _GEN_22151 = io_i_ex_res_packs_0_valid ? _GEN_19975 : _GEN_17798; // @[rob.scala 141:39]
  wire [4:0] _GEN_22152 = io_i_ex_res_packs_0_valid ? _GEN_19976 : _GEN_17799; // @[rob.scala 141:39]
  wire [4:0] _GEN_22153 = io_i_ex_res_packs_0_valid ? _GEN_19977 : _GEN_17800; // @[rob.scala 141:39]
  wire [4:0] _GEN_22154 = io_i_ex_res_packs_0_valid ? _GEN_19978 : _GEN_17801; // @[rob.scala 141:39]
  wire [4:0] _GEN_22155 = io_i_ex_res_packs_0_valid ? _GEN_19979 : _GEN_17802; // @[rob.scala 141:39]
  wire [4:0] _GEN_22156 = io_i_ex_res_packs_0_valid ? _GEN_19980 : _GEN_17803; // @[rob.scala 141:39]
  wire [4:0] _GEN_22157 = io_i_ex_res_packs_0_valid ? _GEN_19981 : _GEN_17804; // @[rob.scala 141:39]
  wire [4:0] _GEN_22158 = io_i_ex_res_packs_0_valid ? _GEN_19982 : _GEN_17805; // @[rob.scala 141:39]
  wire [4:0] _GEN_22159 = io_i_ex_res_packs_0_valid ? _GEN_19983 : _GEN_17806; // @[rob.scala 141:39]
  wire [4:0] _GEN_22160 = io_i_ex_res_packs_0_valid ? _GEN_19984 : _GEN_17807; // @[rob.scala 141:39]
  wire [4:0] _GEN_22161 = io_i_ex_res_packs_0_valid ? _GEN_19985 : _GEN_17808; // @[rob.scala 141:39]
  wire [4:0] _GEN_22162 = io_i_ex_res_packs_0_valid ? _GEN_19986 : _GEN_17809; // @[rob.scala 141:39]
  wire [4:0] _GEN_22163 = io_i_ex_res_packs_0_valid ? _GEN_19987 : _GEN_17810; // @[rob.scala 141:39]
  wire [4:0] _GEN_22164 = io_i_ex_res_packs_0_valid ? _GEN_19988 : _GEN_17811; // @[rob.scala 141:39]
  wire [4:0] _GEN_22165 = io_i_ex_res_packs_0_valid ? _GEN_19989 : _GEN_17812; // @[rob.scala 141:39]
  wire [4:0] _GEN_22166 = io_i_ex_res_packs_0_valid ? _GEN_19990 : _GEN_17813; // @[rob.scala 141:39]
  wire [4:0] _GEN_22167 = io_i_ex_res_packs_0_valid ? _GEN_19991 : _GEN_17814; // @[rob.scala 141:39]
  wire [4:0] _GEN_22168 = io_i_ex_res_packs_0_valid ? _GEN_19992 : _GEN_17815; // @[rob.scala 141:39]
  wire [4:0] _GEN_22169 = io_i_ex_res_packs_0_valid ? _GEN_19993 : _GEN_17816; // @[rob.scala 141:39]
  wire [4:0] _GEN_22170 = io_i_ex_res_packs_0_valid ? _GEN_19994 : _GEN_17817; // @[rob.scala 141:39]
  wire [4:0] _GEN_22171 = io_i_ex_res_packs_0_valid ? _GEN_19995 : _GEN_17818; // @[rob.scala 141:39]
  wire [4:0] _GEN_22172 = io_i_ex_res_packs_0_valid ? _GEN_19996 : _GEN_17819; // @[rob.scala 141:39]
  wire [4:0] _GEN_22173 = io_i_ex_res_packs_0_valid ? _GEN_19997 : _GEN_17820; // @[rob.scala 141:39]
  wire [4:0] _GEN_22174 = io_i_ex_res_packs_0_valid ? _GEN_19998 : _GEN_17821; // @[rob.scala 141:39]
  wire [4:0] _GEN_22175 = io_i_ex_res_packs_0_valid ? _GEN_19999 : _GEN_17822; // @[rob.scala 141:39]
  wire [4:0] _GEN_22176 = io_i_ex_res_packs_0_valid ? _GEN_20000 : _GEN_17823; // @[rob.scala 141:39]
  wire [4:0] _GEN_22177 = io_i_ex_res_packs_0_valid ? _GEN_20001 : _GEN_17824; // @[rob.scala 141:39]
  wire [4:0] _GEN_22178 = io_i_ex_res_packs_0_valid ? _GEN_20002 : _GEN_17825; // @[rob.scala 141:39]
  wire [4:0] _GEN_22179 = io_i_ex_res_packs_0_valid ? _GEN_20003 : _GEN_17826; // @[rob.scala 141:39]
  wire [4:0] _GEN_22180 = io_i_ex_res_packs_0_valid ? _GEN_20004 : _GEN_17827; // @[rob.scala 141:39]
  wire [4:0] _GEN_22181 = io_i_ex_res_packs_0_valid ? _GEN_20005 : _GEN_17828; // @[rob.scala 141:39]
  wire [4:0] _GEN_22182 = io_i_ex_res_packs_0_valid ? _GEN_20006 : _GEN_17829; // @[rob.scala 141:39]
  wire [4:0] _GEN_22183 = io_i_ex_res_packs_0_valid ? _GEN_20007 : _GEN_17830; // @[rob.scala 141:39]
  wire [4:0] _GEN_22184 = io_i_ex_res_packs_0_valid ? _GEN_20008 : _GEN_17831; // @[rob.scala 141:39]
  wire [4:0] _GEN_22185 = io_i_ex_res_packs_0_valid ? _GEN_20009 : _GEN_17832; // @[rob.scala 141:39]
  wire [4:0] _GEN_22186 = io_i_ex_res_packs_0_valid ? _GEN_20010 : _GEN_17833; // @[rob.scala 141:39]
  wire [4:0] _GEN_22187 = io_i_ex_res_packs_0_valid ? _GEN_20011 : _GEN_17834; // @[rob.scala 141:39]
  wire [4:0] _GEN_22188 = io_i_ex_res_packs_0_valid ? _GEN_20012 : _GEN_17835; // @[rob.scala 141:39]
  wire [4:0] _GEN_22189 = io_i_ex_res_packs_0_valid ? _GEN_20013 : _GEN_17836; // @[rob.scala 141:39]
  wire [4:0] _GEN_22190 = io_i_ex_res_packs_0_valid ? _GEN_20014 : _GEN_17837; // @[rob.scala 141:39]
  wire [4:0] _GEN_22191 = io_i_ex_res_packs_0_valid ? _GEN_20015 : _GEN_17838; // @[rob.scala 141:39]
  wire [4:0] _GEN_22192 = io_i_ex_res_packs_0_valid ? _GEN_20016 : _GEN_17839; // @[rob.scala 141:39]
  wire [4:0] _GEN_22193 = io_i_ex_res_packs_0_valid ? _GEN_20017 : _GEN_17840; // @[rob.scala 141:39]
  wire [4:0] _GEN_22194 = io_i_ex_res_packs_0_valid ? _GEN_20018 : _GEN_17841; // @[rob.scala 141:39]
  wire [4:0] _GEN_22195 = io_i_ex_res_packs_0_valid ? _GEN_20019 : _GEN_17842; // @[rob.scala 141:39]
  wire [4:0] _GEN_22196 = io_i_ex_res_packs_0_valid ? _GEN_20020 : _GEN_17843; // @[rob.scala 141:39]
  wire [4:0] _GEN_22197 = io_i_ex_res_packs_0_valid ? _GEN_20021 : _GEN_17844; // @[rob.scala 141:39]
  wire [4:0] _GEN_22198 = io_i_ex_res_packs_0_valid ? _GEN_20022 : _GEN_17845; // @[rob.scala 141:39]
  wire [4:0] _GEN_22199 = io_i_ex_res_packs_0_valid ? _GEN_20023 : _GEN_17846; // @[rob.scala 141:39]
  wire [4:0] _GEN_22200 = io_i_ex_res_packs_0_valid ? _GEN_20024 : _GEN_17847; // @[rob.scala 141:39]
  wire [4:0] _GEN_22201 = io_i_ex_res_packs_0_valid ? _GEN_20025 : _GEN_17848; // @[rob.scala 141:39]
  wire [4:0] _GEN_22202 = io_i_ex_res_packs_0_valid ? _GEN_20026 : _GEN_17849; // @[rob.scala 141:39]
  wire [4:0] _GEN_22203 = io_i_ex_res_packs_0_valid ? _GEN_20027 : _GEN_17850; // @[rob.scala 141:39]
  wire [4:0] _GEN_22204 = io_i_ex_res_packs_0_valid ? _GEN_20028 : _GEN_17851; // @[rob.scala 141:39]
  wire [4:0] _GEN_22205 = io_i_ex_res_packs_0_valid ? _GEN_20029 : _GEN_17852; // @[rob.scala 141:39]
  wire [4:0] _GEN_22206 = io_i_ex_res_packs_0_valid ? _GEN_20030 : _GEN_17853; // @[rob.scala 141:39]
  wire [4:0] _GEN_22207 = io_i_ex_res_packs_0_valid ? _GEN_20031 : _GEN_17854; // @[rob.scala 141:39]
  wire [4:0] _GEN_22208 = io_i_ex_res_packs_0_valid ? _GEN_20032 : _GEN_17855; // @[rob.scala 141:39]
  wire [4:0] _GEN_22209 = io_i_ex_res_packs_0_valid ? _GEN_20033 : _GEN_17856; // @[rob.scala 141:39]
  wire [63:0] _GEN_22850 = io_i_ex_res_packs_0_valid ? _GEN_20674 : _GEN_18497; // @[rob.scala 141:39]
  wire [63:0] _GEN_22851 = io_i_ex_res_packs_0_valid ? _GEN_20675 : _GEN_18498; // @[rob.scala 141:39]
  wire [63:0] _GEN_22852 = io_i_ex_res_packs_0_valid ? _GEN_20676 : _GEN_18499; // @[rob.scala 141:39]
  wire [63:0] _GEN_22853 = io_i_ex_res_packs_0_valid ? _GEN_20677 : _GEN_18500; // @[rob.scala 141:39]
  wire [63:0] _GEN_22854 = io_i_ex_res_packs_0_valid ? _GEN_20678 : _GEN_18501; // @[rob.scala 141:39]
  wire [63:0] _GEN_22855 = io_i_ex_res_packs_0_valid ? _GEN_20679 : _GEN_18502; // @[rob.scala 141:39]
  wire [63:0] _GEN_22856 = io_i_ex_res_packs_0_valid ? _GEN_20680 : _GEN_18503; // @[rob.scala 141:39]
  wire [63:0] _GEN_22857 = io_i_ex_res_packs_0_valid ? _GEN_20681 : _GEN_18504; // @[rob.scala 141:39]
  wire [63:0] _GEN_22858 = io_i_ex_res_packs_0_valid ? _GEN_20682 : _GEN_18505; // @[rob.scala 141:39]
  wire [63:0] _GEN_22859 = io_i_ex_res_packs_0_valid ? _GEN_20683 : _GEN_18506; // @[rob.scala 141:39]
  wire [63:0] _GEN_22860 = io_i_ex_res_packs_0_valid ? _GEN_20684 : _GEN_18507; // @[rob.scala 141:39]
  wire [63:0] _GEN_22861 = io_i_ex_res_packs_0_valid ? _GEN_20685 : _GEN_18508; // @[rob.scala 141:39]
  wire [63:0] _GEN_22862 = io_i_ex_res_packs_0_valid ? _GEN_20686 : _GEN_18509; // @[rob.scala 141:39]
  wire [63:0] _GEN_22863 = io_i_ex_res_packs_0_valid ? _GEN_20687 : _GEN_18510; // @[rob.scala 141:39]
  wire [63:0] _GEN_22864 = io_i_ex_res_packs_0_valid ? _GEN_20688 : _GEN_18511; // @[rob.scala 141:39]
  wire [63:0] _GEN_22865 = io_i_ex_res_packs_0_valid ? _GEN_20689 : _GEN_18512; // @[rob.scala 141:39]
  wire [63:0] _GEN_22866 = io_i_ex_res_packs_0_valid ? _GEN_20690 : _GEN_18513; // @[rob.scala 141:39]
  wire [63:0] _GEN_22867 = io_i_ex_res_packs_0_valid ? _GEN_20691 : _GEN_18514; // @[rob.scala 141:39]
  wire [63:0] _GEN_22868 = io_i_ex_res_packs_0_valid ? _GEN_20692 : _GEN_18515; // @[rob.scala 141:39]
  wire [63:0] _GEN_22869 = io_i_ex_res_packs_0_valid ? _GEN_20693 : _GEN_18516; // @[rob.scala 141:39]
  wire [63:0] _GEN_22870 = io_i_ex_res_packs_0_valid ? _GEN_20694 : _GEN_18517; // @[rob.scala 141:39]
  wire [63:0] _GEN_22871 = io_i_ex_res_packs_0_valid ? _GEN_20695 : _GEN_18518; // @[rob.scala 141:39]
  wire [63:0] _GEN_22872 = io_i_ex_res_packs_0_valid ? _GEN_20696 : _GEN_18519; // @[rob.scala 141:39]
  wire [63:0] _GEN_22873 = io_i_ex_res_packs_0_valid ? _GEN_20697 : _GEN_18520; // @[rob.scala 141:39]
  wire [63:0] _GEN_22874 = io_i_ex_res_packs_0_valid ? _GEN_20698 : _GEN_18521; // @[rob.scala 141:39]
  wire [63:0] _GEN_22875 = io_i_ex_res_packs_0_valid ? _GEN_20699 : _GEN_18522; // @[rob.scala 141:39]
  wire [63:0] _GEN_22876 = io_i_ex_res_packs_0_valid ? _GEN_20700 : _GEN_18523; // @[rob.scala 141:39]
  wire [63:0] _GEN_22877 = io_i_ex_res_packs_0_valid ? _GEN_20701 : _GEN_18524; // @[rob.scala 141:39]
  wire [63:0] _GEN_22878 = io_i_ex_res_packs_0_valid ? _GEN_20702 : _GEN_18525; // @[rob.scala 141:39]
  wire [63:0] _GEN_22879 = io_i_ex_res_packs_0_valid ? _GEN_20703 : _GEN_18526; // @[rob.scala 141:39]
  wire [63:0] _GEN_22880 = io_i_ex_res_packs_0_valid ? _GEN_20704 : _GEN_18527; // @[rob.scala 141:39]
  wire [63:0] _GEN_22881 = io_i_ex_res_packs_0_valid ? _GEN_20705 : _GEN_18528; // @[rob.scala 141:39]
  wire [63:0] _GEN_22882 = io_i_ex_res_packs_0_valid ? _GEN_20706 : _GEN_18529; // @[rob.scala 141:39]
  wire [63:0] _GEN_22883 = io_i_ex_res_packs_0_valid ? _GEN_20707 : _GEN_18530; // @[rob.scala 141:39]
  wire [63:0] _GEN_22884 = io_i_ex_res_packs_0_valid ? _GEN_20708 : _GEN_18531; // @[rob.scala 141:39]
  wire [63:0] _GEN_22885 = io_i_ex_res_packs_0_valid ? _GEN_20709 : _GEN_18532; // @[rob.scala 141:39]
  wire [63:0] _GEN_22886 = io_i_ex_res_packs_0_valid ? _GEN_20710 : _GEN_18533; // @[rob.scala 141:39]
  wire [63:0] _GEN_22887 = io_i_ex_res_packs_0_valid ? _GEN_20711 : _GEN_18534; // @[rob.scala 141:39]
  wire [63:0] _GEN_22888 = io_i_ex_res_packs_0_valid ? _GEN_20712 : _GEN_18535; // @[rob.scala 141:39]
  wire [63:0] _GEN_22889 = io_i_ex_res_packs_0_valid ? _GEN_20713 : _GEN_18536; // @[rob.scala 141:39]
  wire [63:0] _GEN_22890 = io_i_ex_res_packs_0_valid ? _GEN_20714 : _GEN_18537; // @[rob.scala 141:39]
  wire [63:0] _GEN_22891 = io_i_ex_res_packs_0_valid ? _GEN_20715 : _GEN_18538; // @[rob.scala 141:39]
  wire [63:0] _GEN_22892 = io_i_ex_res_packs_0_valid ? _GEN_20716 : _GEN_18539; // @[rob.scala 141:39]
  wire [63:0] _GEN_22893 = io_i_ex_res_packs_0_valid ? _GEN_20717 : _GEN_18540; // @[rob.scala 141:39]
  wire [63:0] _GEN_22894 = io_i_ex_res_packs_0_valid ? _GEN_20718 : _GEN_18541; // @[rob.scala 141:39]
  wire [63:0] _GEN_22895 = io_i_ex_res_packs_0_valid ? _GEN_20719 : _GEN_18542; // @[rob.scala 141:39]
  wire [63:0] _GEN_22896 = io_i_ex_res_packs_0_valid ? _GEN_20720 : _GEN_18543; // @[rob.scala 141:39]
  wire [63:0] _GEN_22897 = io_i_ex_res_packs_0_valid ? _GEN_20721 : _GEN_18544; // @[rob.scala 141:39]
  wire [63:0] _GEN_22898 = io_i_ex_res_packs_0_valid ? _GEN_20722 : _GEN_18545; // @[rob.scala 141:39]
  wire [63:0] _GEN_22899 = io_i_ex_res_packs_0_valid ? _GEN_20723 : _GEN_18546; // @[rob.scala 141:39]
  wire [63:0] _GEN_22900 = io_i_ex_res_packs_0_valid ? _GEN_20724 : _GEN_18547; // @[rob.scala 141:39]
  wire [63:0] _GEN_22901 = io_i_ex_res_packs_0_valid ? _GEN_20725 : _GEN_18548; // @[rob.scala 141:39]
  wire [63:0] _GEN_22902 = io_i_ex_res_packs_0_valid ? _GEN_20726 : _GEN_18549; // @[rob.scala 141:39]
  wire [63:0] _GEN_22903 = io_i_ex_res_packs_0_valid ? _GEN_20727 : _GEN_18550; // @[rob.scala 141:39]
  wire [63:0] _GEN_22904 = io_i_ex_res_packs_0_valid ? _GEN_20728 : _GEN_18551; // @[rob.scala 141:39]
  wire [63:0] _GEN_22905 = io_i_ex_res_packs_0_valid ? _GEN_20729 : _GEN_18552; // @[rob.scala 141:39]
  wire [63:0] _GEN_22906 = io_i_ex_res_packs_0_valid ? _GEN_20730 : _GEN_18553; // @[rob.scala 141:39]
  wire [63:0] _GEN_22907 = io_i_ex_res_packs_0_valid ? _GEN_20731 : _GEN_18554; // @[rob.scala 141:39]
  wire [63:0] _GEN_22908 = io_i_ex_res_packs_0_valid ? _GEN_20732 : _GEN_18555; // @[rob.scala 141:39]
  wire [63:0] _GEN_22909 = io_i_ex_res_packs_0_valid ? _GEN_20733 : _GEN_18556; // @[rob.scala 141:39]
  wire [63:0] _GEN_22910 = io_i_ex_res_packs_0_valid ? _GEN_20734 : _GEN_18557; // @[rob.scala 141:39]
  wire [63:0] _GEN_22911 = io_i_ex_res_packs_0_valid ? _GEN_20735 : _GEN_18558; // @[rob.scala 141:39]
  wire [63:0] _GEN_22912 = io_i_ex_res_packs_0_valid ? _GEN_20736 : _GEN_18559; // @[rob.scala 141:39]
  wire [63:0] _GEN_22913 = io_i_ex_res_packs_0_valid ? _GEN_20737 : _GEN_18560; // @[rob.scala 141:39]
  wire [63:0] _GEN_22914 = io_i_ex_res_packs_0_valid ? _GEN_20738 : _GEN_18561; // @[rob.scala 141:39]
  wire [63:0] _GEN_22915 = io_i_ex_res_packs_0_valid ? _GEN_20739 : _GEN_18562; // @[rob.scala 141:39]
  wire [63:0] _GEN_22916 = io_i_ex_res_packs_0_valid ? _GEN_20740 : _GEN_18563; // @[rob.scala 141:39]
  wire [63:0] _GEN_22917 = io_i_ex_res_packs_0_valid ? _GEN_20741 : _GEN_18564; // @[rob.scala 141:39]
  wire [63:0] _GEN_22918 = io_i_ex_res_packs_0_valid ? _GEN_20742 : _GEN_18565; // @[rob.scala 141:39]
  wire [63:0] _GEN_22919 = io_i_ex_res_packs_0_valid ? _GEN_20743 : _GEN_18566; // @[rob.scala 141:39]
  wire [63:0] _GEN_22920 = io_i_ex_res_packs_0_valid ? _GEN_20744 : _GEN_18567; // @[rob.scala 141:39]
  wire [63:0] _GEN_22921 = io_i_ex_res_packs_0_valid ? _GEN_20745 : _GEN_18568; // @[rob.scala 141:39]
  wire [63:0] _GEN_22922 = io_i_ex_res_packs_0_valid ? _GEN_20746 : _GEN_18569; // @[rob.scala 141:39]
  wire [63:0] _GEN_22923 = io_i_ex_res_packs_0_valid ? _GEN_20747 : _GEN_18570; // @[rob.scala 141:39]
  wire [63:0] _GEN_22924 = io_i_ex_res_packs_0_valid ? _GEN_20748 : _GEN_18571; // @[rob.scala 141:39]
  wire [63:0] _GEN_22925 = io_i_ex_res_packs_0_valid ? _GEN_20749 : _GEN_18572; // @[rob.scala 141:39]
  wire [63:0] _GEN_22926 = io_i_ex_res_packs_0_valid ? _GEN_20750 : _GEN_18573; // @[rob.scala 141:39]
  wire [63:0] _GEN_22927 = io_i_ex_res_packs_0_valid ? _GEN_20751 : _GEN_18574; // @[rob.scala 141:39]
  wire [63:0] _GEN_22928 = io_i_ex_res_packs_0_valid ? _GEN_20752 : _GEN_18575; // @[rob.scala 141:39]
  wire [63:0] _GEN_22929 = io_i_ex_res_packs_0_valid ? _GEN_20753 : _GEN_18576; // @[rob.scala 141:39]
  wire [63:0] _GEN_22930 = io_i_ex_res_packs_0_valid ? _GEN_20754 : _GEN_18577; // @[rob.scala 141:39]
  wire [63:0] _GEN_22931 = io_i_ex_res_packs_0_valid ? _GEN_20755 : _GEN_18578; // @[rob.scala 141:39]
  wire [63:0] _GEN_22932 = io_i_ex_res_packs_0_valid ? _GEN_20756 : _GEN_18579; // @[rob.scala 141:39]
  wire [63:0] _GEN_22933 = io_i_ex_res_packs_0_valid ? _GEN_20757 : _GEN_18580; // @[rob.scala 141:39]
  wire [63:0] _GEN_22934 = io_i_ex_res_packs_0_valid ? _GEN_20758 : _GEN_18581; // @[rob.scala 141:39]
  wire [63:0] _GEN_22935 = io_i_ex_res_packs_0_valid ? _GEN_20759 : _GEN_18582; // @[rob.scala 141:39]
  wire [63:0] _GEN_22936 = io_i_ex_res_packs_0_valid ? _GEN_20760 : _GEN_18583; // @[rob.scala 141:39]
  wire [63:0] _GEN_22937 = io_i_ex_res_packs_0_valid ? _GEN_20761 : _GEN_18584; // @[rob.scala 141:39]
  wire [63:0] _GEN_22938 = io_i_ex_res_packs_0_valid ? _GEN_20762 : _GEN_18585; // @[rob.scala 141:39]
  wire [63:0] _GEN_22939 = io_i_ex_res_packs_0_valid ? _GEN_20763 : _GEN_18586; // @[rob.scala 141:39]
  wire [63:0] _GEN_22940 = io_i_ex_res_packs_0_valid ? _GEN_20764 : _GEN_18587; // @[rob.scala 141:39]
  wire [63:0] _GEN_22941 = io_i_ex_res_packs_0_valid ? _GEN_20765 : _GEN_18588; // @[rob.scala 141:39]
  wire [63:0] _GEN_22942 = io_i_ex_res_packs_0_valid ? _GEN_20766 : _GEN_18589; // @[rob.scala 141:39]
  wire [63:0] _GEN_22943 = io_i_ex_res_packs_0_valid ? _GEN_20767 : _GEN_18590; // @[rob.scala 141:39]
  wire [63:0] _GEN_22944 = io_i_ex_res_packs_0_valid ? _GEN_20768 : _GEN_18591; // @[rob.scala 141:39]
  wire [63:0] _GEN_22945 = io_i_ex_res_packs_0_valid ? _GEN_20769 : _GEN_18592; // @[rob.scala 141:39]
  wire [63:0] _GEN_22946 = io_i_ex_res_packs_0_valid ? _GEN_20770 : _GEN_18593; // @[rob.scala 141:39]
  wire [63:0] _GEN_22947 = io_i_ex_res_packs_0_valid ? _GEN_20771 : _GEN_18594; // @[rob.scala 141:39]
  wire [63:0] _GEN_22948 = io_i_ex_res_packs_0_valid ? _GEN_20772 : _GEN_18595; // @[rob.scala 141:39]
  wire [63:0] _GEN_22949 = io_i_ex_res_packs_0_valid ? _GEN_20773 : _GEN_18596; // @[rob.scala 141:39]
  wire [63:0] _GEN_22950 = io_i_ex_res_packs_0_valid ? _GEN_20774 : _GEN_18597; // @[rob.scala 141:39]
  wire [63:0] _GEN_22951 = io_i_ex_res_packs_0_valid ? _GEN_20775 : _GEN_18598; // @[rob.scala 141:39]
  wire [63:0] _GEN_22952 = io_i_ex_res_packs_0_valid ? _GEN_20776 : _GEN_18599; // @[rob.scala 141:39]
  wire [63:0] _GEN_22953 = io_i_ex_res_packs_0_valid ? _GEN_20777 : _GEN_18600; // @[rob.scala 141:39]
  wire [63:0] _GEN_22954 = io_i_ex_res_packs_0_valid ? _GEN_20778 : _GEN_18601; // @[rob.scala 141:39]
  wire [63:0] _GEN_22955 = io_i_ex_res_packs_0_valid ? _GEN_20779 : _GEN_18602; // @[rob.scala 141:39]
  wire [63:0] _GEN_22956 = io_i_ex_res_packs_0_valid ? _GEN_20780 : _GEN_18603; // @[rob.scala 141:39]
  wire [63:0] _GEN_22957 = io_i_ex_res_packs_0_valid ? _GEN_20781 : _GEN_18604; // @[rob.scala 141:39]
  wire [63:0] _GEN_22958 = io_i_ex_res_packs_0_valid ? _GEN_20782 : _GEN_18605; // @[rob.scala 141:39]
  wire [63:0] _GEN_22959 = io_i_ex_res_packs_0_valid ? _GEN_20783 : _GEN_18606; // @[rob.scala 141:39]
  wire [63:0] _GEN_22960 = io_i_ex_res_packs_0_valid ? _GEN_20784 : _GEN_18607; // @[rob.scala 141:39]
  wire [63:0] _GEN_22961 = io_i_ex_res_packs_0_valid ? _GEN_20785 : _GEN_18608; // @[rob.scala 141:39]
  wire [63:0] _GEN_22962 = io_i_ex_res_packs_0_valid ? _GEN_20786 : _GEN_18609; // @[rob.scala 141:39]
  wire [63:0] _GEN_22963 = io_i_ex_res_packs_0_valid ? _GEN_20787 : _GEN_18610; // @[rob.scala 141:39]
  wire [63:0] _GEN_22964 = io_i_ex_res_packs_0_valid ? _GEN_20788 : _GEN_18611; // @[rob.scala 141:39]
  wire [63:0] _GEN_22965 = io_i_ex_res_packs_0_valid ? _GEN_20789 : _GEN_18612; // @[rob.scala 141:39]
  wire [63:0] _GEN_22966 = io_i_ex_res_packs_0_valid ? _GEN_20790 : _GEN_18613; // @[rob.scala 141:39]
  wire [63:0] _GEN_22967 = io_i_ex_res_packs_0_valid ? _GEN_20791 : _GEN_18614; // @[rob.scala 141:39]
  wire [63:0] _GEN_22968 = io_i_ex_res_packs_0_valid ? _GEN_20792 : _GEN_18615; // @[rob.scala 141:39]
  wire [63:0] _GEN_22969 = io_i_ex_res_packs_0_valid ? _GEN_20793 : _GEN_18616; // @[rob.scala 141:39]
  wire [63:0] _GEN_22970 = io_i_ex_res_packs_0_valid ? _GEN_20794 : _GEN_18617; // @[rob.scala 141:39]
  wire [63:0] _GEN_22971 = io_i_ex_res_packs_0_valid ? _GEN_20795 : _GEN_18618; // @[rob.scala 141:39]
  wire [63:0] _GEN_22972 = io_i_ex_res_packs_0_valid ? _GEN_20796 : _GEN_18619; // @[rob.scala 141:39]
  wire [63:0] _GEN_22973 = io_i_ex_res_packs_0_valid ? _GEN_20797 : _GEN_18620; // @[rob.scala 141:39]
  wire [63:0] _GEN_22974 = io_i_ex_res_packs_0_valid ? _GEN_20798 : _GEN_18621; // @[rob.scala 141:39]
  wire [63:0] _GEN_22975 = io_i_ex_res_packs_0_valid ? _GEN_20799 : _GEN_18622; // @[rob.scala 141:39]
  wire [63:0] _GEN_22976 = io_i_ex_res_packs_0_valid ? _GEN_20800 : _GEN_18623; // @[rob.scala 141:39]
  wire [63:0] _GEN_22977 = io_i_ex_res_packs_0_valid ? _GEN_20801 : _GEN_18624; // @[rob.scala 141:39]
  wire [4:0] _GEN_23234 = io_i_ex_res_packs_0_valid ? _GEN_21058 : _GEN_18881; // @[rob.scala 141:39]
  wire [4:0] _GEN_23235 = io_i_ex_res_packs_0_valid ? _GEN_21059 : _GEN_18882; // @[rob.scala 141:39]
  wire [4:0] _GEN_23236 = io_i_ex_res_packs_0_valid ? _GEN_21060 : _GEN_18883; // @[rob.scala 141:39]
  wire [4:0] _GEN_23237 = io_i_ex_res_packs_0_valid ? _GEN_21061 : _GEN_18884; // @[rob.scala 141:39]
  wire [4:0] _GEN_23238 = io_i_ex_res_packs_0_valid ? _GEN_21062 : _GEN_18885; // @[rob.scala 141:39]
  wire [4:0] _GEN_23239 = io_i_ex_res_packs_0_valid ? _GEN_21063 : _GEN_18886; // @[rob.scala 141:39]
  wire [4:0] _GEN_23240 = io_i_ex_res_packs_0_valid ? _GEN_21064 : _GEN_18887; // @[rob.scala 141:39]
  wire [4:0] _GEN_23241 = io_i_ex_res_packs_0_valid ? _GEN_21065 : _GEN_18888; // @[rob.scala 141:39]
  wire [4:0] _GEN_23242 = io_i_ex_res_packs_0_valid ? _GEN_21066 : _GEN_18889; // @[rob.scala 141:39]
  wire [4:0] _GEN_23243 = io_i_ex_res_packs_0_valid ? _GEN_21067 : _GEN_18890; // @[rob.scala 141:39]
  wire [4:0] _GEN_23244 = io_i_ex_res_packs_0_valid ? _GEN_21068 : _GEN_18891; // @[rob.scala 141:39]
  wire [4:0] _GEN_23245 = io_i_ex_res_packs_0_valid ? _GEN_21069 : _GEN_18892; // @[rob.scala 141:39]
  wire [4:0] _GEN_23246 = io_i_ex_res_packs_0_valid ? _GEN_21070 : _GEN_18893; // @[rob.scala 141:39]
  wire [4:0] _GEN_23247 = io_i_ex_res_packs_0_valid ? _GEN_21071 : _GEN_18894; // @[rob.scala 141:39]
  wire [4:0] _GEN_23248 = io_i_ex_res_packs_0_valid ? _GEN_21072 : _GEN_18895; // @[rob.scala 141:39]
  wire [4:0] _GEN_23249 = io_i_ex_res_packs_0_valid ? _GEN_21073 : _GEN_18896; // @[rob.scala 141:39]
  wire [4:0] _GEN_23250 = io_i_ex_res_packs_0_valid ? _GEN_21074 : _GEN_18897; // @[rob.scala 141:39]
  wire [4:0] _GEN_23251 = io_i_ex_res_packs_0_valid ? _GEN_21075 : _GEN_18898; // @[rob.scala 141:39]
  wire [4:0] _GEN_23252 = io_i_ex_res_packs_0_valid ? _GEN_21076 : _GEN_18899; // @[rob.scala 141:39]
  wire [4:0] _GEN_23253 = io_i_ex_res_packs_0_valid ? _GEN_21077 : _GEN_18900; // @[rob.scala 141:39]
  wire [4:0] _GEN_23254 = io_i_ex_res_packs_0_valid ? _GEN_21078 : _GEN_18901; // @[rob.scala 141:39]
  wire [4:0] _GEN_23255 = io_i_ex_res_packs_0_valid ? _GEN_21079 : _GEN_18902; // @[rob.scala 141:39]
  wire [4:0] _GEN_23256 = io_i_ex_res_packs_0_valid ? _GEN_21080 : _GEN_18903; // @[rob.scala 141:39]
  wire [4:0] _GEN_23257 = io_i_ex_res_packs_0_valid ? _GEN_21081 : _GEN_18904; // @[rob.scala 141:39]
  wire [4:0] _GEN_23258 = io_i_ex_res_packs_0_valid ? _GEN_21082 : _GEN_18905; // @[rob.scala 141:39]
  wire [4:0] _GEN_23259 = io_i_ex_res_packs_0_valid ? _GEN_21083 : _GEN_18906; // @[rob.scala 141:39]
  wire [4:0] _GEN_23260 = io_i_ex_res_packs_0_valid ? _GEN_21084 : _GEN_18907; // @[rob.scala 141:39]
  wire [4:0] _GEN_23261 = io_i_ex_res_packs_0_valid ? _GEN_21085 : _GEN_18908; // @[rob.scala 141:39]
  wire [4:0] _GEN_23262 = io_i_ex_res_packs_0_valid ? _GEN_21086 : _GEN_18909; // @[rob.scala 141:39]
  wire [4:0] _GEN_23263 = io_i_ex_res_packs_0_valid ? _GEN_21087 : _GEN_18910; // @[rob.scala 141:39]
  wire [4:0] _GEN_23264 = io_i_ex_res_packs_0_valid ? _GEN_21088 : _GEN_18911; // @[rob.scala 141:39]
  wire [4:0] _GEN_23265 = io_i_ex_res_packs_0_valid ? _GEN_21089 : _GEN_18912; // @[rob.scala 141:39]
  wire [4:0] _GEN_23266 = io_i_ex_res_packs_0_valid ? _GEN_21090 : _GEN_18913; // @[rob.scala 141:39]
  wire [4:0] _GEN_23267 = io_i_ex_res_packs_0_valid ? _GEN_21091 : _GEN_18914; // @[rob.scala 141:39]
  wire [4:0] _GEN_23268 = io_i_ex_res_packs_0_valid ? _GEN_21092 : _GEN_18915; // @[rob.scala 141:39]
  wire [4:0] _GEN_23269 = io_i_ex_res_packs_0_valid ? _GEN_21093 : _GEN_18916; // @[rob.scala 141:39]
  wire [4:0] _GEN_23270 = io_i_ex_res_packs_0_valid ? _GEN_21094 : _GEN_18917; // @[rob.scala 141:39]
  wire [4:0] _GEN_23271 = io_i_ex_res_packs_0_valid ? _GEN_21095 : _GEN_18918; // @[rob.scala 141:39]
  wire [4:0] _GEN_23272 = io_i_ex_res_packs_0_valid ? _GEN_21096 : _GEN_18919; // @[rob.scala 141:39]
  wire [4:0] _GEN_23273 = io_i_ex_res_packs_0_valid ? _GEN_21097 : _GEN_18920; // @[rob.scala 141:39]
  wire [4:0] _GEN_23274 = io_i_ex_res_packs_0_valid ? _GEN_21098 : _GEN_18921; // @[rob.scala 141:39]
  wire [4:0] _GEN_23275 = io_i_ex_res_packs_0_valid ? _GEN_21099 : _GEN_18922; // @[rob.scala 141:39]
  wire [4:0] _GEN_23276 = io_i_ex_res_packs_0_valid ? _GEN_21100 : _GEN_18923; // @[rob.scala 141:39]
  wire [4:0] _GEN_23277 = io_i_ex_res_packs_0_valid ? _GEN_21101 : _GEN_18924; // @[rob.scala 141:39]
  wire [4:0] _GEN_23278 = io_i_ex_res_packs_0_valid ? _GEN_21102 : _GEN_18925; // @[rob.scala 141:39]
  wire [4:0] _GEN_23279 = io_i_ex_res_packs_0_valid ? _GEN_21103 : _GEN_18926; // @[rob.scala 141:39]
  wire [4:0] _GEN_23280 = io_i_ex_res_packs_0_valid ? _GEN_21104 : _GEN_18927; // @[rob.scala 141:39]
  wire [4:0] _GEN_23281 = io_i_ex_res_packs_0_valid ? _GEN_21105 : _GEN_18928; // @[rob.scala 141:39]
  wire [4:0] _GEN_23282 = io_i_ex_res_packs_0_valid ? _GEN_21106 : _GEN_18929; // @[rob.scala 141:39]
  wire [4:0] _GEN_23283 = io_i_ex_res_packs_0_valid ? _GEN_21107 : _GEN_18930; // @[rob.scala 141:39]
  wire [4:0] _GEN_23284 = io_i_ex_res_packs_0_valid ? _GEN_21108 : _GEN_18931; // @[rob.scala 141:39]
  wire [4:0] _GEN_23285 = io_i_ex_res_packs_0_valid ? _GEN_21109 : _GEN_18932; // @[rob.scala 141:39]
  wire [4:0] _GEN_23286 = io_i_ex_res_packs_0_valid ? _GEN_21110 : _GEN_18933; // @[rob.scala 141:39]
  wire [4:0] _GEN_23287 = io_i_ex_res_packs_0_valid ? _GEN_21111 : _GEN_18934; // @[rob.scala 141:39]
  wire [4:0] _GEN_23288 = io_i_ex_res_packs_0_valid ? _GEN_21112 : _GEN_18935; // @[rob.scala 141:39]
  wire [4:0] _GEN_23289 = io_i_ex_res_packs_0_valid ? _GEN_21113 : _GEN_18936; // @[rob.scala 141:39]
  wire [4:0] _GEN_23290 = io_i_ex_res_packs_0_valid ? _GEN_21114 : _GEN_18937; // @[rob.scala 141:39]
  wire [4:0] _GEN_23291 = io_i_ex_res_packs_0_valid ? _GEN_21115 : _GEN_18938; // @[rob.scala 141:39]
  wire [4:0] _GEN_23292 = io_i_ex_res_packs_0_valid ? _GEN_21116 : _GEN_18939; // @[rob.scala 141:39]
  wire [4:0] _GEN_23293 = io_i_ex_res_packs_0_valid ? _GEN_21117 : _GEN_18940; // @[rob.scala 141:39]
  wire [4:0] _GEN_23294 = io_i_ex_res_packs_0_valid ? _GEN_21118 : _GEN_18941; // @[rob.scala 141:39]
  wire [4:0] _GEN_23295 = io_i_ex_res_packs_0_valid ? _GEN_21119 : _GEN_18942; // @[rob.scala 141:39]
  wire [4:0] _GEN_23296 = io_i_ex_res_packs_0_valid ? _GEN_21120 : _GEN_18943; // @[rob.scala 141:39]
  wire [4:0] _GEN_23297 = io_i_ex_res_packs_0_valid ? _GEN_21121 : _GEN_18944; // @[rob.scala 141:39]
  wire  _GEN_23490 = io_i_ex_res_packs_0_valid ? _GEN_21314 : _GEN_19137; // @[rob.scala 141:39]
  wire  _GEN_23491 = io_i_ex_res_packs_0_valid ? _GEN_21315 : _GEN_19138; // @[rob.scala 141:39]
  wire  _GEN_23492 = io_i_ex_res_packs_0_valid ? _GEN_21316 : _GEN_19139; // @[rob.scala 141:39]
  wire  _GEN_23493 = io_i_ex_res_packs_0_valid ? _GEN_21317 : _GEN_19140; // @[rob.scala 141:39]
  wire  _GEN_23494 = io_i_ex_res_packs_0_valid ? _GEN_21318 : _GEN_19141; // @[rob.scala 141:39]
  wire  _GEN_23495 = io_i_ex_res_packs_0_valid ? _GEN_21319 : _GEN_19142; // @[rob.scala 141:39]
  wire  _GEN_23496 = io_i_ex_res_packs_0_valid ? _GEN_21320 : _GEN_19143; // @[rob.scala 141:39]
  wire  _GEN_23497 = io_i_ex_res_packs_0_valid ? _GEN_21321 : _GEN_19144; // @[rob.scala 141:39]
  wire  _GEN_23498 = io_i_ex_res_packs_0_valid ? _GEN_21322 : _GEN_19145; // @[rob.scala 141:39]
  wire  _GEN_23499 = io_i_ex_res_packs_0_valid ? _GEN_21323 : _GEN_19146; // @[rob.scala 141:39]
  wire  _GEN_23500 = io_i_ex_res_packs_0_valid ? _GEN_21324 : _GEN_19147; // @[rob.scala 141:39]
  wire  _GEN_23501 = io_i_ex_res_packs_0_valid ? _GEN_21325 : _GEN_19148; // @[rob.scala 141:39]
  wire  _GEN_23502 = io_i_ex_res_packs_0_valid ? _GEN_21326 : _GEN_19149; // @[rob.scala 141:39]
  wire  _GEN_23503 = io_i_ex_res_packs_0_valid ? _GEN_21327 : _GEN_19150; // @[rob.scala 141:39]
  wire  _GEN_23504 = io_i_ex_res_packs_0_valid ? _GEN_21328 : _GEN_19151; // @[rob.scala 141:39]
  wire  _GEN_23505 = io_i_ex_res_packs_0_valid ? _GEN_21329 : _GEN_19152; // @[rob.scala 141:39]
  wire  _GEN_23506 = io_i_ex_res_packs_0_valid ? _GEN_21330 : _GEN_19153; // @[rob.scala 141:39]
  wire  _GEN_23507 = io_i_ex_res_packs_0_valid ? _GEN_21331 : _GEN_19154; // @[rob.scala 141:39]
  wire  _GEN_23508 = io_i_ex_res_packs_0_valid ? _GEN_21332 : _GEN_19155; // @[rob.scala 141:39]
  wire  _GEN_23509 = io_i_ex_res_packs_0_valid ? _GEN_21333 : _GEN_19156; // @[rob.scala 141:39]
  wire  _GEN_23510 = io_i_ex_res_packs_0_valid ? _GEN_21334 : _GEN_19157; // @[rob.scala 141:39]
  wire  _GEN_23511 = io_i_ex_res_packs_0_valid ? _GEN_21335 : _GEN_19158; // @[rob.scala 141:39]
  wire  _GEN_23512 = io_i_ex_res_packs_0_valid ? _GEN_21336 : _GEN_19159; // @[rob.scala 141:39]
  wire  _GEN_23513 = io_i_ex_res_packs_0_valid ? _GEN_21337 : _GEN_19160; // @[rob.scala 141:39]
  wire  _GEN_23514 = io_i_ex_res_packs_0_valid ? _GEN_21338 : _GEN_19161; // @[rob.scala 141:39]
  wire  _GEN_23515 = io_i_ex_res_packs_0_valid ? _GEN_21339 : _GEN_19162; // @[rob.scala 141:39]
  wire  _GEN_23516 = io_i_ex_res_packs_0_valid ? _GEN_21340 : _GEN_19163; // @[rob.scala 141:39]
  wire  _GEN_23517 = io_i_ex_res_packs_0_valid ? _GEN_21341 : _GEN_19164; // @[rob.scala 141:39]
  wire  _GEN_23518 = io_i_ex_res_packs_0_valid ? _GEN_21342 : _GEN_19165; // @[rob.scala 141:39]
  wire  _GEN_23519 = io_i_ex_res_packs_0_valid ? _GEN_21343 : _GEN_19166; // @[rob.scala 141:39]
  wire  _GEN_23520 = io_i_ex_res_packs_0_valid ? _GEN_21344 : _GEN_19167; // @[rob.scala 141:39]
  wire  _GEN_23521 = io_i_ex_res_packs_0_valid ? _GEN_21345 : _GEN_19168; // @[rob.scala 141:39]
  wire  _GEN_23522 = io_i_ex_res_packs_0_valid ? _GEN_21346 : _GEN_19169; // @[rob.scala 141:39]
  wire  _GEN_23523 = io_i_ex_res_packs_0_valid ? _GEN_21347 : _GEN_19170; // @[rob.scala 141:39]
  wire  _GEN_23524 = io_i_ex_res_packs_0_valid ? _GEN_21348 : _GEN_19171; // @[rob.scala 141:39]
  wire  _GEN_23525 = io_i_ex_res_packs_0_valid ? _GEN_21349 : _GEN_19172; // @[rob.scala 141:39]
  wire  _GEN_23526 = io_i_ex_res_packs_0_valid ? _GEN_21350 : _GEN_19173; // @[rob.scala 141:39]
  wire  _GEN_23527 = io_i_ex_res_packs_0_valid ? _GEN_21351 : _GEN_19174; // @[rob.scala 141:39]
  wire  _GEN_23528 = io_i_ex_res_packs_0_valid ? _GEN_21352 : _GEN_19175; // @[rob.scala 141:39]
  wire  _GEN_23529 = io_i_ex_res_packs_0_valid ? _GEN_21353 : _GEN_19176; // @[rob.scala 141:39]
  wire  _GEN_23530 = io_i_ex_res_packs_0_valid ? _GEN_21354 : _GEN_19177; // @[rob.scala 141:39]
  wire  _GEN_23531 = io_i_ex_res_packs_0_valid ? _GEN_21355 : _GEN_19178; // @[rob.scala 141:39]
  wire  _GEN_23532 = io_i_ex_res_packs_0_valid ? _GEN_21356 : _GEN_19179; // @[rob.scala 141:39]
  wire  _GEN_23533 = io_i_ex_res_packs_0_valid ? _GEN_21357 : _GEN_19180; // @[rob.scala 141:39]
  wire  _GEN_23534 = io_i_ex_res_packs_0_valid ? _GEN_21358 : _GEN_19181; // @[rob.scala 141:39]
  wire  _GEN_23535 = io_i_ex_res_packs_0_valid ? _GEN_21359 : _GEN_19182; // @[rob.scala 141:39]
  wire  _GEN_23536 = io_i_ex_res_packs_0_valid ? _GEN_21360 : _GEN_19183; // @[rob.scala 141:39]
  wire  _GEN_23537 = io_i_ex_res_packs_0_valid ? _GEN_21361 : _GEN_19184; // @[rob.scala 141:39]
  wire  _GEN_23538 = io_i_ex_res_packs_0_valid ? _GEN_21362 : _GEN_19185; // @[rob.scala 141:39]
  wire  _GEN_23539 = io_i_ex_res_packs_0_valid ? _GEN_21363 : _GEN_19186; // @[rob.scala 141:39]
  wire  _GEN_23540 = io_i_ex_res_packs_0_valid ? _GEN_21364 : _GEN_19187; // @[rob.scala 141:39]
  wire  _GEN_23541 = io_i_ex_res_packs_0_valid ? _GEN_21365 : _GEN_19188; // @[rob.scala 141:39]
  wire  _GEN_23542 = io_i_ex_res_packs_0_valid ? _GEN_21366 : _GEN_19189; // @[rob.scala 141:39]
  wire  _GEN_23543 = io_i_ex_res_packs_0_valid ? _GEN_21367 : _GEN_19190; // @[rob.scala 141:39]
  wire  _GEN_23544 = io_i_ex_res_packs_0_valid ? _GEN_21368 : _GEN_19191; // @[rob.scala 141:39]
  wire  _GEN_23545 = io_i_ex_res_packs_0_valid ? _GEN_21369 : _GEN_19192; // @[rob.scala 141:39]
  wire  _GEN_23546 = io_i_ex_res_packs_0_valid ? _GEN_21370 : _GEN_19193; // @[rob.scala 141:39]
  wire  _GEN_23547 = io_i_ex_res_packs_0_valid ? _GEN_21371 : _GEN_19194; // @[rob.scala 141:39]
  wire  _GEN_23548 = io_i_ex_res_packs_0_valid ? _GEN_21372 : _GEN_19195; // @[rob.scala 141:39]
  wire  _GEN_23549 = io_i_ex_res_packs_0_valid ? _GEN_21373 : _GEN_19196; // @[rob.scala 141:39]
  wire  _GEN_23550 = io_i_ex_res_packs_0_valid ? _GEN_21374 : _GEN_19197; // @[rob.scala 141:39]
  wire  _GEN_23551 = io_i_ex_res_packs_0_valid ? _GEN_21375 : _GEN_19198; // @[rob.scala 141:39]
  wire  _GEN_23552 = io_i_ex_res_packs_0_valid ? _GEN_21376 : _GEN_19199; // @[rob.scala 141:39]
  wire  _GEN_23553 = io_i_ex_res_packs_0_valid ? _GEN_21377 : _GEN_19200; // @[rob.scala 141:39]
  wire  _GEN_42193 = 6'h0 == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23554 = 6'h0 == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21378; // @[rob.scala 148:{53,53}]
  wire  _GEN_42194 = 6'h1 == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23555 = 6'h1 == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21379; // @[rob.scala 148:{53,53}]
  wire  _GEN_42195 = 6'h2 == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23556 = 6'h2 == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21380; // @[rob.scala 148:{53,53}]
  wire  _GEN_42196 = 6'h3 == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23557 = 6'h3 == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21381; // @[rob.scala 148:{53,53}]
  wire  _GEN_42197 = 6'h4 == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23558 = 6'h4 == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21382; // @[rob.scala 148:{53,53}]
  wire  _GEN_42198 = 6'h5 == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23559 = 6'h5 == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21383; // @[rob.scala 148:{53,53}]
  wire  _GEN_42199 = 6'h6 == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23560 = 6'h6 == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21384; // @[rob.scala 148:{53,53}]
  wire  _GEN_42200 = 6'h7 == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23561 = 6'h7 == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21385; // @[rob.scala 148:{53,53}]
  wire  _GEN_42201 = 6'h8 == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23562 = 6'h8 == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21386; // @[rob.scala 148:{53,53}]
  wire  _GEN_42202 = 6'h9 == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23563 = 6'h9 == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21387; // @[rob.scala 148:{53,53}]
  wire  _GEN_42203 = 6'ha == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23564 = 6'ha == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21388; // @[rob.scala 148:{53,53}]
  wire  _GEN_42204 = 6'hb == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23565 = 6'hb == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21389; // @[rob.scala 148:{53,53}]
  wire  _GEN_42205 = 6'hc == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23566 = 6'hc == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21390; // @[rob.scala 148:{53,53}]
  wire  _GEN_42206 = 6'hd == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23567 = 6'hd == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21391; // @[rob.scala 148:{53,53}]
  wire  _GEN_42207 = 6'he == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23568 = 6'he == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21392; // @[rob.scala 148:{53,53}]
  wire  _GEN_42208 = 6'hf == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23569 = 6'hf == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21393; // @[rob.scala 148:{53,53}]
  wire  _GEN_42209 = 6'h10 == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23570 = 6'h10 == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21394; // @[rob.scala 148:{53,53}]
  wire  _GEN_42210 = 6'h11 == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23571 = 6'h11 == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21395; // @[rob.scala 148:{53,53}]
  wire  _GEN_42211 = 6'h12 == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23572 = 6'h12 == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21396; // @[rob.scala 148:{53,53}]
  wire  _GEN_42212 = 6'h13 == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23573 = 6'h13 == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21397; // @[rob.scala 148:{53,53}]
  wire  _GEN_42213 = 6'h14 == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23574 = 6'h14 == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21398; // @[rob.scala 148:{53,53}]
  wire  _GEN_42214 = 6'h15 == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23575 = 6'h15 == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21399; // @[rob.scala 148:{53,53}]
  wire  _GEN_42215 = 6'h16 == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23576 = 6'h16 == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21400; // @[rob.scala 148:{53,53}]
  wire  _GEN_42216 = 6'h17 == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23577 = 6'h17 == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21401; // @[rob.scala 148:{53,53}]
  wire  _GEN_42217 = 6'h18 == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23578 = 6'h18 == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21402; // @[rob.scala 148:{53,53}]
  wire  _GEN_42218 = 6'h19 == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23579 = 6'h19 == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21403; // @[rob.scala 148:{53,53}]
  wire  _GEN_42219 = 6'h1a == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23580 = 6'h1a == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21404; // @[rob.scala 148:{53,53}]
  wire  _GEN_42220 = 6'h1b == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23581 = 6'h1b == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21405; // @[rob.scala 148:{53,53}]
  wire  _GEN_42221 = 6'h1c == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23582 = 6'h1c == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21406; // @[rob.scala 148:{53,53}]
  wire  _GEN_42222 = 6'h1d == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23583 = 6'h1d == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21407; // @[rob.scala 148:{53,53}]
  wire  _GEN_42223 = 6'h1e == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23584 = 6'h1e == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21408; // @[rob.scala 148:{53,53}]
  wire  _GEN_42224 = 6'h1f == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23585 = 6'h1f == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21409; // @[rob.scala 148:{53,53}]
  wire  _GEN_42225 = 6'h20 == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23586 = 6'h20 == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21410; // @[rob.scala 148:{53,53}]
  wire  _GEN_42226 = 6'h21 == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23587 = 6'h21 == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21411; // @[rob.scala 148:{53,53}]
  wire  _GEN_42227 = 6'h22 == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23588 = 6'h22 == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21412; // @[rob.scala 148:{53,53}]
  wire  _GEN_42228 = 6'h23 == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23589 = 6'h23 == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21413; // @[rob.scala 148:{53,53}]
  wire  _GEN_42229 = 6'h24 == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23590 = 6'h24 == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21414; // @[rob.scala 148:{53,53}]
  wire  _GEN_42230 = 6'h25 == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23591 = 6'h25 == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21415; // @[rob.scala 148:{53,53}]
  wire  _GEN_42231 = 6'h26 == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23592 = 6'h26 == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21416; // @[rob.scala 148:{53,53}]
  wire  _GEN_42232 = 6'h27 == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23593 = 6'h27 == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21417; // @[rob.scala 148:{53,53}]
  wire  _GEN_42233 = 6'h28 == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23594 = 6'h28 == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21418; // @[rob.scala 148:{53,53}]
  wire  _GEN_42234 = 6'h29 == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23595 = 6'h29 == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21419; // @[rob.scala 148:{53,53}]
  wire  _GEN_42235 = 6'h2a == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23596 = 6'h2a == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21420; // @[rob.scala 148:{53,53}]
  wire  _GEN_42236 = 6'h2b == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23597 = 6'h2b == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21421; // @[rob.scala 148:{53,53}]
  wire  _GEN_42237 = 6'h2c == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23598 = 6'h2c == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21422; // @[rob.scala 148:{53,53}]
  wire  _GEN_42238 = 6'h2d == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23599 = 6'h2d == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21423; // @[rob.scala 148:{53,53}]
  wire  _GEN_42239 = 6'h2e == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23600 = 6'h2e == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21424; // @[rob.scala 148:{53,53}]
  wire  _GEN_42240 = 6'h2f == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23601 = 6'h2f == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21425; // @[rob.scala 148:{53,53}]
  wire  _GEN_42241 = 6'h30 == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23602 = 6'h30 == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21426; // @[rob.scala 148:{53,53}]
  wire  _GEN_42242 = 6'h31 == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23603 = 6'h31 == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21427; // @[rob.scala 148:{53,53}]
  wire  _GEN_42243 = 6'h32 == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23604 = 6'h32 == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21428; // @[rob.scala 148:{53,53}]
  wire  _GEN_42244 = 6'h33 == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23605 = 6'h33 == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21429; // @[rob.scala 148:{53,53}]
  wire  _GEN_42245 = 6'h34 == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23606 = 6'h34 == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21430; // @[rob.scala 148:{53,53}]
  wire  _GEN_42246 = 6'h35 == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23607 = 6'h35 == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21431; // @[rob.scala 148:{53,53}]
  wire  _GEN_42247 = 6'h36 == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23608 = 6'h36 == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21432; // @[rob.scala 148:{53,53}]
  wire  _GEN_42248 = 6'h37 == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23609 = 6'h37 == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21433; // @[rob.scala 148:{53,53}]
  wire  _GEN_42249 = 6'h38 == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23610 = 6'h38 == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21434; // @[rob.scala 148:{53,53}]
  wire  _GEN_42250 = 6'h39 == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23611 = 6'h39 == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21435; // @[rob.scala 148:{53,53}]
  wire  _GEN_42251 = 6'h3a == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23612 = 6'h3a == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21436; // @[rob.scala 148:{53,53}]
  wire  _GEN_42252 = 6'h3b == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23613 = 6'h3b == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21437; // @[rob.scala 148:{53,53}]
  wire  _GEN_42253 = 6'h3c == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23614 = 6'h3c == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21438; // @[rob.scala 148:{53,53}]
  wire  _GEN_42254 = 6'h3d == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23615 = 6'h3d == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21439; // @[rob.scala 148:{53,53}]
  wire  _GEN_42255 = 6'h3e == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23616 = 6'h3e == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21440; // @[rob.scala 148:{53,53}]
  wire  _GEN_42256 = 6'h3f == io_i_ex_res_packs_1_uop_rob_idx[5:0]; // @[rob.scala 148:{53,53}]
  wire  _GEN_23617 = 6'h3f == io_i_ex_res_packs_1_uop_rob_idx[5:0] | _GEN_21441; // @[rob.scala 148:{53,53}]
  wire [31:0] _GEN_23682 = 6'h0 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21506; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23683 = 6'h1 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21507; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23684 = 6'h2 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21508; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23685 = 6'h3 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21509; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23686 = 6'h4 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21510; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23687 = 6'h5 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21511; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23688 = 6'h6 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21512; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23689 = 6'h7 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21513; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23690 = 6'h8 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21514; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23691 = 6'h9 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21515; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23692 = 6'ha == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21516; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23693 = 6'hb == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21517; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23694 = 6'hc == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21518; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23695 = 6'hd == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21519; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23696 = 6'he == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21520; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23697 = 6'hf == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21521; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23698 = 6'h10 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21522; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23699 = 6'h11 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21523; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23700 = 6'h12 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21524; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23701 = 6'h13 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21525; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23702 = 6'h14 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21526; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23703 = 6'h15 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21527; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23704 = 6'h16 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21528; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23705 = 6'h17 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21529; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23706 = 6'h18 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21530; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23707 = 6'h19 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21531; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23708 = 6'h1a == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21532; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23709 = 6'h1b == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21533; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23710 = 6'h1c == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21534; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23711 = 6'h1d == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21535; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23712 = 6'h1e == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21536; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23713 = 6'h1f == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21537; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23714 = 6'h20 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21538; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23715 = 6'h21 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21539; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23716 = 6'h22 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21540; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23717 = 6'h23 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21541; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23718 = 6'h24 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21542; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23719 = 6'h25 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21543; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23720 = 6'h26 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21544; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23721 = 6'h27 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21545; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23722 = 6'h28 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21546; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23723 = 6'h29 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21547; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23724 = 6'h2a == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21548; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23725 = 6'h2b == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21549; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23726 = 6'h2c == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21550; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23727 = 6'h2d == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21551; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23728 = 6'h2e == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21552; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23729 = 6'h2f == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21553; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23730 = 6'h30 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21554; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23731 = 6'h31 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21555; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23732 = 6'h32 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21556; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23733 = 6'h33 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21557; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23734 = 6'h34 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21558; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23735 = 6'h35 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21559; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23736 = 6'h36 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21560; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23737 = 6'h37 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21561; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23738 = 6'h38 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21562; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23739 = 6'h39 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21563; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23740 = 6'h3a == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21564; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23741 = 6'h3b == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21565; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23742 = 6'h3c == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21566; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23743 = 6'h3d == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21567; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23744 = 6'h3e == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21568; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23745 = 6'h3f == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_pc : _GEN_21569; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23746 = 6'h0 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21570; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23747 = 6'h1 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21571; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23748 = 6'h2 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21572; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23749 = 6'h3 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21573; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23750 = 6'h4 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21574; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23751 = 6'h5 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21575; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23752 = 6'h6 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21576; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23753 = 6'h7 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21577; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23754 = 6'h8 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21578; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23755 = 6'h9 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21579; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23756 = 6'ha == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21580; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23757 = 6'hb == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21581; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23758 = 6'hc == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21582; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23759 = 6'hd == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21583; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23760 = 6'he == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21584; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23761 = 6'hf == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21585; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23762 = 6'h10 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21586; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23763 = 6'h11 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21587; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23764 = 6'h12 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21588; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23765 = 6'h13 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21589; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23766 = 6'h14 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21590; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23767 = 6'h15 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21591; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23768 = 6'h16 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21592; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23769 = 6'h17 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21593; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23770 = 6'h18 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21594; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23771 = 6'h19 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21595; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23772 = 6'h1a == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21596; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23773 = 6'h1b == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21597; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23774 = 6'h1c == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21598; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23775 = 6'h1d == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21599; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23776 = 6'h1e == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21600; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23777 = 6'h1f == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21601; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23778 = 6'h20 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21602; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23779 = 6'h21 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21603; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23780 = 6'h22 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21604; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23781 = 6'h23 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21605; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23782 = 6'h24 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21606; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23783 = 6'h25 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21607; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23784 = 6'h26 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21608; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23785 = 6'h27 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21609; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23786 = 6'h28 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21610; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23787 = 6'h29 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21611; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23788 = 6'h2a == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21612; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23789 = 6'h2b == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21613; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23790 = 6'h2c == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21614; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23791 = 6'h2d == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21615; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23792 = 6'h2e == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21616; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23793 = 6'h2f == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21617; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23794 = 6'h30 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21618; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23795 = 6'h31 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21619; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23796 = 6'h32 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21620; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23797 = 6'h33 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21621; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23798 = 6'h34 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21622; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23799 = 6'h35 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21623; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23800 = 6'h36 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21624; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23801 = 6'h37 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21625; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23802 = 6'h38 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21626; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23803 = 6'h39 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21627; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23804 = 6'h3a == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21628; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23805 = 6'h3b == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21629; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23806 = 6'h3c == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21630; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23807 = 6'h3d == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21631; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23808 = 6'h3e == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21632; // @[rob.scala 149:{51,51}]
  wire [31:0] _GEN_23809 = 6'h3f == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_inst : _GEN_21633; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23810 = 6'h0 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21634; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23811 = 6'h1 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21635; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23812 = 6'h2 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21636; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23813 = 6'h3 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21637; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23814 = 6'h4 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21638; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23815 = 6'h5 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21639; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23816 = 6'h6 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21640; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23817 = 6'h7 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21641; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23818 = 6'h8 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21642; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23819 = 6'h9 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21643; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23820 = 6'ha == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21644; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23821 = 6'hb == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21645; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23822 = 6'hc == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21646; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23823 = 6'hd == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21647; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23824 = 6'he == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21648; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23825 = 6'hf == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21649; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23826 = 6'h10 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21650
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23827 = 6'h11 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21651
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23828 = 6'h12 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21652
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23829 = 6'h13 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21653
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23830 = 6'h14 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21654
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23831 = 6'h15 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21655
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23832 = 6'h16 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21656
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23833 = 6'h17 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21657
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23834 = 6'h18 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21658
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23835 = 6'h19 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21659
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23836 = 6'h1a == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21660
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23837 = 6'h1b == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21661
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23838 = 6'h1c == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21662
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23839 = 6'h1d == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21663
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23840 = 6'h1e == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21664
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23841 = 6'h1f == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21665
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23842 = 6'h20 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21666
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23843 = 6'h21 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21667
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23844 = 6'h22 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21668
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23845 = 6'h23 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21669
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23846 = 6'h24 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21670
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23847 = 6'h25 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21671
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23848 = 6'h26 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21672
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23849 = 6'h27 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21673
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23850 = 6'h28 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21674
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23851 = 6'h29 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21675
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23852 = 6'h2a == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21676
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23853 = 6'h2b == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21677
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23854 = 6'h2c == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21678
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23855 = 6'h2d == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21679
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23856 = 6'h2e == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21680
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23857 = 6'h2f == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21681
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23858 = 6'h30 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21682
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23859 = 6'h31 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21683
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23860 = 6'h32 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21684
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23861 = 6'h33 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21685
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23862 = 6'h34 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21686
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23863 = 6'h35 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21687
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23864 = 6'h36 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21688
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23865 = 6'h37 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21689
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23866 = 6'h38 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21690
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23867 = 6'h39 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21691
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23868 = 6'h3a == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21692
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23869 = 6'h3b == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21693
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23870 = 6'h3c == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21694
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23871 = 6'h3d == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21695
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23872 = 6'h3e == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21696
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_23873 = 6'h3f == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_func_code : _GEN_21697
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24194 = 6'h0 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22018; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24195 = 6'h1 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22019; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24196 = 6'h2 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22020; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24197 = 6'h3 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22021; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24198 = 6'h4 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22022; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24199 = 6'h5 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22023; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24200 = 6'h6 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22024; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24201 = 6'h7 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22025; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24202 = 6'h8 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22026; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24203 = 6'h9 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22027; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24204 = 6'ha == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22028; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24205 = 6'hb == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22029; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24206 = 6'hc == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22030; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24207 = 6'hd == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22031; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24208 = 6'he == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22032; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24209 = 6'hf == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22033; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24210 = 6'h10 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22034; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24211 = 6'h11 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22035; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24212 = 6'h12 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22036; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24213 = 6'h13 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22037; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24214 = 6'h14 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22038; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24215 = 6'h15 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22039; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24216 = 6'h16 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22040; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24217 = 6'h17 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22041; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24218 = 6'h18 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22042; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24219 = 6'h19 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22043; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24220 = 6'h1a == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22044; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24221 = 6'h1b == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22045; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24222 = 6'h1c == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22046; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24223 = 6'h1d == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22047; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24224 = 6'h1e == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22048; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24225 = 6'h1f == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22049; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24226 = 6'h20 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22050; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24227 = 6'h21 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22051; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24228 = 6'h22 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22052; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24229 = 6'h23 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22053; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24230 = 6'h24 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22054; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24231 = 6'h25 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22055; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24232 = 6'h26 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22056; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24233 = 6'h27 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22057; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24234 = 6'h28 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22058; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24235 = 6'h29 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22059; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24236 = 6'h2a == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22060; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24237 = 6'h2b == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22061; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24238 = 6'h2c == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22062; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24239 = 6'h2d == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22063; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24240 = 6'h2e == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22064; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24241 = 6'h2f == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22065; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24242 = 6'h30 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22066; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24243 = 6'h31 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22067; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24244 = 6'h32 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22068; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24245 = 6'h33 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22069; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24246 = 6'h34 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22070; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24247 = 6'h35 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22071; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24248 = 6'h36 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22072; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24249 = 6'h37 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22073; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24250 = 6'h38 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22074; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24251 = 6'h39 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22075; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24252 = 6'h3a == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22076; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24253 = 6'h3b == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22077; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24254 = 6'h3c == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22078; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24255 = 6'h3d == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22079; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24256 = 6'h3e == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22080; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24257 = 6'h3f == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_phy_dst : _GEN_22081; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24258 = 6'h0 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22082; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24259 = 6'h1 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22083; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24260 = 6'h2 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22084; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24261 = 6'h3 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22085; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24262 = 6'h4 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22086; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24263 = 6'h5 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22087; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24264 = 6'h6 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22088; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24265 = 6'h7 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22089; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24266 = 6'h8 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22090; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24267 = 6'h9 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22091; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24268 = 6'ha == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22092; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24269 = 6'hb == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22093; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24270 = 6'hc == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22094; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24271 = 6'hd == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22095; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24272 = 6'he == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22096; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24273 = 6'hf == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22097; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24274 = 6'h10 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22098
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24275 = 6'h11 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22099
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24276 = 6'h12 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22100
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24277 = 6'h13 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22101
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24278 = 6'h14 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22102
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24279 = 6'h15 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22103
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24280 = 6'h16 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22104
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24281 = 6'h17 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22105
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24282 = 6'h18 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22106
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24283 = 6'h19 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22107
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24284 = 6'h1a == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22108
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24285 = 6'h1b == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22109
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24286 = 6'h1c == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22110
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24287 = 6'h1d == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22111
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24288 = 6'h1e == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22112
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24289 = 6'h1f == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22113
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24290 = 6'h20 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22114
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24291 = 6'h21 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22115
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24292 = 6'h22 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22116
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24293 = 6'h23 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22117
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24294 = 6'h24 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22118
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24295 = 6'h25 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22119
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24296 = 6'h26 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22120
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24297 = 6'h27 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22121
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24298 = 6'h28 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22122
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24299 = 6'h29 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22123
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24300 = 6'h2a == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22124
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24301 = 6'h2b == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22125
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24302 = 6'h2c == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22126
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24303 = 6'h2d == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22127
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24304 = 6'h2e == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22128
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24305 = 6'h2f == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22129
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24306 = 6'h30 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22130
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24307 = 6'h31 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22131
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24308 = 6'h32 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22132
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24309 = 6'h33 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22133
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24310 = 6'h34 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22134
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24311 = 6'h35 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22135
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24312 = 6'h36 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22136
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24313 = 6'h37 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22137
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24314 = 6'h38 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22138
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24315 = 6'h39 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22139
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24316 = 6'h3a == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22140
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24317 = 6'h3b == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22141
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24318 = 6'h3c == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22142
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24319 = 6'h3d == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22143
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24320 = 6'h3e == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22144
    ; // @[rob.scala 149:{51,51}]
  wire [6:0] _GEN_24321 = 6'h3f == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_stale_dst : _GEN_22145
    ; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24322 = 6'h0 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22146; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24323 = 6'h1 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22147; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24324 = 6'h2 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22148; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24325 = 6'h3 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22149; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24326 = 6'h4 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22150; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24327 = 6'h5 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22151; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24328 = 6'h6 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22152; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24329 = 6'h7 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22153; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24330 = 6'h8 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22154; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24331 = 6'h9 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22155; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24332 = 6'ha == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22156; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24333 = 6'hb == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22157; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24334 = 6'hc == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22158; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24335 = 6'hd == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22159; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24336 = 6'he == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22160; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24337 = 6'hf == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22161; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24338 = 6'h10 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22162; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24339 = 6'h11 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22163; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24340 = 6'h12 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22164; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24341 = 6'h13 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22165; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24342 = 6'h14 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22166; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24343 = 6'h15 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22167; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24344 = 6'h16 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22168; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24345 = 6'h17 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22169; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24346 = 6'h18 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22170; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24347 = 6'h19 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22171; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24348 = 6'h1a == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22172; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24349 = 6'h1b == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22173; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24350 = 6'h1c == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22174; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24351 = 6'h1d == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22175; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24352 = 6'h1e == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22176; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24353 = 6'h1f == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22177; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24354 = 6'h20 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22178; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24355 = 6'h21 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22179; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24356 = 6'h22 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22180; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24357 = 6'h23 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22181; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24358 = 6'h24 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22182; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24359 = 6'h25 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22183; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24360 = 6'h26 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22184; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24361 = 6'h27 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22185; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24362 = 6'h28 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22186; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24363 = 6'h29 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22187; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24364 = 6'h2a == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22188; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24365 = 6'h2b == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22189; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24366 = 6'h2c == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22190; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24367 = 6'h2d == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22191; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24368 = 6'h2e == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22192; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24369 = 6'h2f == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22193; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24370 = 6'h30 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22194; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24371 = 6'h31 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22195; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24372 = 6'h32 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22196; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24373 = 6'h33 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22197; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24374 = 6'h34 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22198; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24375 = 6'h35 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22199; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24376 = 6'h36 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22200; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24377 = 6'h37 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22201; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24378 = 6'h38 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22202; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24379 = 6'h39 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22203; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24380 = 6'h3a == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22204; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24381 = 6'h3b == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22205; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24382 = 6'h3c == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22206; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24383 = 6'h3d == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22207; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24384 = 6'h3e == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22208; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_24385 = 6'h3f == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_arch_dst : _GEN_22209; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25026 = 6'h0 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value : _GEN_22850
    ; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25027 = 6'h1 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value : _GEN_22851
    ; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25028 = 6'h2 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value : _GEN_22852
    ; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25029 = 6'h3 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value : _GEN_22853
    ; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25030 = 6'h4 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value : _GEN_22854
    ; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25031 = 6'h5 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value : _GEN_22855
    ; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25032 = 6'h6 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value : _GEN_22856
    ; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25033 = 6'h7 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value : _GEN_22857
    ; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25034 = 6'h8 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value : _GEN_22858
    ; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25035 = 6'h9 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value : _GEN_22859
    ; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25036 = 6'ha == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value : _GEN_22860
    ; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25037 = 6'hb == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value : _GEN_22861
    ; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25038 = 6'hc == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value : _GEN_22862
    ; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25039 = 6'hd == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value : _GEN_22863
    ; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25040 = 6'he == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value : _GEN_22864
    ; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25041 = 6'hf == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value : _GEN_22865
    ; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25042 = 6'h10 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22866; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25043 = 6'h11 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22867; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25044 = 6'h12 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22868; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25045 = 6'h13 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22869; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25046 = 6'h14 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22870; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25047 = 6'h15 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22871; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25048 = 6'h16 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22872; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25049 = 6'h17 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22873; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25050 = 6'h18 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22874; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25051 = 6'h19 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22875; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25052 = 6'h1a == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22876; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25053 = 6'h1b == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22877; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25054 = 6'h1c == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22878; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25055 = 6'h1d == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22879; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25056 = 6'h1e == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22880; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25057 = 6'h1f == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22881; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25058 = 6'h20 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22882; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25059 = 6'h21 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22883; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25060 = 6'h22 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22884; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25061 = 6'h23 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22885; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25062 = 6'h24 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22886; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25063 = 6'h25 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22887; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25064 = 6'h26 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22888; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25065 = 6'h27 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22889; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25066 = 6'h28 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22890; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25067 = 6'h29 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22891; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25068 = 6'h2a == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22892; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25069 = 6'h2b == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22893; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25070 = 6'h2c == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22894; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25071 = 6'h2d == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22895; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25072 = 6'h2e == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22896; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25073 = 6'h2f == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22897; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25074 = 6'h30 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22898; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25075 = 6'h31 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22899; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25076 = 6'h32 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22900; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25077 = 6'h33 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22901; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25078 = 6'h34 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22902; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25079 = 6'h35 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22903; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25080 = 6'h36 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22904; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25081 = 6'h37 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22905; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25082 = 6'h38 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22906; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25083 = 6'h39 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22907; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25084 = 6'h3a == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22908; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25085 = 6'h3b == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22909; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25086 = 6'h3c == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22910; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25087 = 6'h3d == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22911; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25088 = 6'h3e == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22912; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25089 = 6'h3f == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_dst_value :
    _GEN_22913; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25090 = 6'h0 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22914; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25091 = 6'h1 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22915; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25092 = 6'h2 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22916; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25093 = 6'h3 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22917; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25094 = 6'h4 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22918; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25095 = 6'h5 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22919; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25096 = 6'h6 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22920; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25097 = 6'h7 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22921; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25098 = 6'h8 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22922; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25099 = 6'h9 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22923; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25100 = 6'ha == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22924; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25101 = 6'hb == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22925; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25102 = 6'hc == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22926; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25103 = 6'hd == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22927; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25104 = 6'he == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22928; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25105 = 6'hf == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22929; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25106 = 6'h10 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22930; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25107 = 6'h11 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22931; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25108 = 6'h12 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22932; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25109 = 6'h13 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22933; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25110 = 6'h14 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22934; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25111 = 6'h15 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22935; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25112 = 6'h16 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22936; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25113 = 6'h17 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22937; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25114 = 6'h18 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22938; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25115 = 6'h19 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22939; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25116 = 6'h1a == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22940; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25117 = 6'h1b == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22941; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25118 = 6'h1c == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22942; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25119 = 6'h1d == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22943; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25120 = 6'h1e == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22944; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25121 = 6'h1f == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22945; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25122 = 6'h20 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22946; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25123 = 6'h21 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22947; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25124 = 6'h22 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22948; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25125 = 6'h23 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22949; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25126 = 6'h24 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22950; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25127 = 6'h25 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22951; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25128 = 6'h26 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22952; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25129 = 6'h27 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22953; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25130 = 6'h28 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22954; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25131 = 6'h29 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22955; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25132 = 6'h2a == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22956; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25133 = 6'h2b == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22957; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25134 = 6'h2c == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22958; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25135 = 6'h2d == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22959; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25136 = 6'h2e == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22960; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25137 = 6'h2f == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22961; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25138 = 6'h30 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22962; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25139 = 6'h31 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22963; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25140 = 6'h32 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22964; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25141 = 6'h33 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22965; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25142 = 6'h34 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22966; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25143 = 6'h35 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22967; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25144 = 6'h36 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22968; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25145 = 6'h37 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22969; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25146 = 6'h38 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22970; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25147 = 6'h39 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22971; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25148 = 6'h3a == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22972; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25149 = 6'h3b == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22973; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25150 = 6'h3c == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22974; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25151 = 6'h3d == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22975; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25152 = 6'h3e == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22976; // @[rob.scala 149:{51,51}]
  wire [63:0] _GEN_25153 = 6'h3f == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_src1_value :
    _GEN_22977; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25410 = 6'h0 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23234; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25411 = 6'h1 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23235; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25412 = 6'h2 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23236; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25413 = 6'h3 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23237; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25414 = 6'h4 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23238; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25415 = 6'h5 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23239; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25416 = 6'h6 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23240; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25417 = 6'h7 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23241; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25418 = 6'h8 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23242; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25419 = 6'h9 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23243; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25420 = 6'ha == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23244; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25421 = 6'hb == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23245; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25422 = 6'hc == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23246; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25423 = 6'hd == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23247; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25424 = 6'he == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23248; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25425 = 6'hf == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23249; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25426 = 6'h10 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23250; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25427 = 6'h11 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23251; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25428 = 6'h12 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23252; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25429 = 6'h13 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23253; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25430 = 6'h14 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23254; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25431 = 6'h15 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23255; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25432 = 6'h16 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23256; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25433 = 6'h17 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23257; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25434 = 6'h18 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23258; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25435 = 6'h19 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23259; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25436 = 6'h1a == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23260; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25437 = 6'h1b == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23261; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25438 = 6'h1c == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23262; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25439 = 6'h1d == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23263; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25440 = 6'h1e == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23264; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25441 = 6'h1f == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23265; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25442 = 6'h20 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23266; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25443 = 6'h21 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23267; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25444 = 6'h22 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23268; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25445 = 6'h23 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23269; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25446 = 6'h24 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23270; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25447 = 6'h25 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23271; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25448 = 6'h26 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23272; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25449 = 6'h27 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23273; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25450 = 6'h28 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23274; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25451 = 6'h29 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23275; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25452 = 6'h2a == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23276; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25453 = 6'h2b == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23277; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25454 = 6'h2c == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23278; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25455 = 6'h2d == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23279; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25456 = 6'h2e == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23280; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25457 = 6'h2f == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23281; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25458 = 6'h30 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23282; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25459 = 6'h31 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23283; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25460 = 6'h32 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23284; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25461 = 6'h33 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23285; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25462 = 6'h34 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23286; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25463 = 6'h35 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23287; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25464 = 6'h36 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23288; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25465 = 6'h37 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23289; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25466 = 6'h38 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23290; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25467 = 6'h39 == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23291; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25468 = 6'h3a == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23292; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25469 = 6'h3b == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23293; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25470 = 6'h3c == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23294; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25471 = 6'h3d == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23295; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25472 = 6'h3e == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23296; // @[rob.scala 149:{51,51}]
  wire [4:0] _GEN_25473 = 6'h3f == io_i_ex_res_packs_1_uop_rob_idx[5:0] ? io_i_ex_res_packs_1_uop_alu_sel : _GEN_23297; // @[rob.scala 149:{51,51}]
  wire  _GEN_25666 = _GEN_42193 | _GEN_23490; // @[rob.scala 151:{52,52}]
  wire  _GEN_25667 = _GEN_42194 | _GEN_23491; // @[rob.scala 151:{52,52}]
  wire  _GEN_25668 = _GEN_42195 | _GEN_23492; // @[rob.scala 151:{52,52}]
  wire  _GEN_25669 = _GEN_42196 | _GEN_23493; // @[rob.scala 151:{52,52}]
  wire  _GEN_25670 = _GEN_42197 | _GEN_23494; // @[rob.scala 151:{52,52}]
  wire  _GEN_25671 = _GEN_42198 | _GEN_23495; // @[rob.scala 151:{52,52}]
  wire  _GEN_25672 = _GEN_42199 | _GEN_23496; // @[rob.scala 151:{52,52}]
  wire  _GEN_25673 = _GEN_42200 | _GEN_23497; // @[rob.scala 151:{52,52}]
  wire  _GEN_25674 = _GEN_42201 | _GEN_23498; // @[rob.scala 151:{52,52}]
  wire  _GEN_25675 = _GEN_42202 | _GEN_23499; // @[rob.scala 151:{52,52}]
  wire  _GEN_25676 = _GEN_42203 | _GEN_23500; // @[rob.scala 151:{52,52}]
  wire  _GEN_25677 = _GEN_42204 | _GEN_23501; // @[rob.scala 151:{52,52}]
  wire  _GEN_25678 = _GEN_42205 | _GEN_23502; // @[rob.scala 151:{52,52}]
  wire  _GEN_25679 = _GEN_42206 | _GEN_23503; // @[rob.scala 151:{52,52}]
  wire  _GEN_25680 = _GEN_42207 | _GEN_23504; // @[rob.scala 151:{52,52}]
  wire  _GEN_25681 = _GEN_42208 | _GEN_23505; // @[rob.scala 151:{52,52}]
  wire  _GEN_25682 = _GEN_42209 | _GEN_23506; // @[rob.scala 151:{52,52}]
  wire  _GEN_25683 = _GEN_42210 | _GEN_23507; // @[rob.scala 151:{52,52}]
  wire  _GEN_25684 = _GEN_42211 | _GEN_23508; // @[rob.scala 151:{52,52}]
  wire  _GEN_25685 = _GEN_42212 | _GEN_23509; // @[rob.scala 151:{52,52}]
  wire  _GEN_25686 = _GEN_42213 | _GEN_23510; // @[rob.scala 151:{52,52}]
  wire  _GEN_25687 = _GEN_42214 | _GEN_23511; // @[rob.scala 151:{52,52}]
  wire  _GEN_25688 = _GEN_42215 | _GEN_23512; // @[rob.scala 151:{52,52}]
  wire  _GEN_25689 = _GEN_42216 | _GEN_23513; // @[rob.scala 151:{52,52}]
  wire  _GEN_25690 = _GEN_42217 | _GEN_23514; // @[rob.scala 151:{52,52}]
  wire  _GEN_25691 = _GEN_42218 | _GEN_23515; // @[rob.scala 151:{52,52}]
  wire  _GEN_25692 = _GEN_42219 | _GEN_23516; // @[rob.scala 151:{52,52}]
  wire  _GEN_25693 = _GEN_42220 | _GEN_23517; // @[rob.scala 151:{52,52}]
  wire  _GEN_25694 = _GEN_42221 | _GEN_23518; // @[rob.scala 151:{52,52}]
  wire  _GEN_25695 = _GEN_42222 | _GEN_23519; // @[rob.scala 151:{52,52}]
  wire  _GEN_25696 = _GEN_42223 | _GEN_23520; // @[rob.scala 151:{52,52}]
  wire  _GEN_25697 = _GEN_42224 | _GEN_23521; // @[rob.scala 151:{52,52}]
  wire  _GEN_25698 = _GEN_42225 | _GEN_23522; // @[rob.scala 151:{52,52}]
  wire  _GEN_25699 = _GEN_42226 | _GEN_23523; // @[rob.scala 151:{52,52}]
  wire  _GEN_25700 = _GEN_42227 | _GEN_23524; // @[rob.scala 151:{52,52}]
  wire  _GEN_25701 = _GEN_42228 | _GEN_23525; // @[rob.scala 151:{52,52}]
  wire  _GEN_25702 = _GEN_42229 | _GEN_23526; // @[rob.scala 151:{52,52}]
  wire  _GEN_25703 = _GEN_42230 | _GEN_23527; // @[rob.scala 151:{52,52}]
  wire  _GEN_25704 = _GEN_42231 | _GEN_23528; // @[rob.scala 151:{52,52}]
  wire  _GEN_25705 = _GEN_42232 | _GEN_23529; // @[rob.scala 151:{52,52}]
  wire  _GEN_25706 = _GEN_42233 | _GEN_23530; // @[rob.scala 151:{52,52}]
  wire  _GEN_25707 = _GEN_42234 | _GEN_23531; // @[rob.scala 151:{52,52}]
  wire  _GEN_25708 = _GEN_42235 | _GEN_23532; // @[rob.scala 151:{52,52}]
  wire  _GEN_25709 = _GEN_42236 | _GEN_23533; // @[rob.scala 151:{52,52}]
  wire  _GEN_25710 = _GEN_42237 | _GEN_23534; // @[rob.scala 151:{52,52}]
  wire  _GEN_25711 = _GEN_42238 | _GEN_23535; // @[rob.scala 151:{52,52}]
  wire  _GEN_25712 = _GEN_42239 | _GEN_23536; // @[rob.scala 151:{52,52}]
  wire  _GEN_25713 = _GEN_42240 | _GEN_23537; // @[rob.scala 151:{52,52}]
  wire  _GEN_25714 = _GEN_42241 | _GEN_23538; // @[rob.scala 151:{52,52}]
  wire  _GEN_25715 = _GEN_42242 | _GEN_23539; // @[rob.scala 151:{52,52}]
  wire  _GEN_25716 = _GEN_42243 | _GEN_23540; // @[rob.scala 151:{52,52}]
  wire  _GEN_25717 = _GEN_42244 | _GEN_23541; // @[rob.scala 151:{52,52}]
  wire  _GEN_25718 = _GEN_42245 | _GEN_23542; // @[rob.scala 151:{52,52}]
  wire  _GEN_25719 = _GEN_42246 | _GEN_23543; // @[rob.scala 151:{52,52}]
  wire  _GEN_25720 = _GEN_42247 | _GEN_23544; // @[rob.scala 151:{52,52}]
  wire  _GEN_25721 = _GEN_42248 | _GEN_23545; // @[rob.scala 151:{52,52}]
  wire  _GEN_25722 = _GEN_42249 | _GEN_23546; // @[rob.scala 151:{52,52}]
  wire  _GEN_25723 = _GEN_42250 | _GEN_23547; // @[rob.scala 151:{52,52}]
  wire  _GEN_25724 = _GEN_42251 | _GEN_23548; // @[rob.scala 151:{52,52}]
  wire  _GEN_25725 = _GEN_42252 | _GEN_23549; // @[rob.scala 151:{52,52}]
  wire  _GEN_25726 = _GEN_42253 | _GEN_23550; // @[rob.scala 151:{52,52}]
  wire  _GEN_25727 = _GEN_42254 | _GEN_23551; // @[rob.scala 151:{52,52}]
  wire  _GEN_25728 = _GEN_42255 | _GEN_23552; // @[rob.scala 151:{52,52}]
  wire  _GEN_25729 = _GEN_42256 | _GEN_23553; // @[rob.scala 151:{52,52}]
  wire  _GEN_25730 = io_i_ex_res_packs_1_valid ? _GEN_23554 : _GEN_21378; // @[rob.scala 147:39]
  wire  _GEN_25731 = io_i_ex_res_packs_1_valid ? _GEN_23555 : _GEN_21379; // @[rob.scala 147:39]
  wire  _GEN_25732 = io_i_ex_res_packs_1_valid ? _GEN_23556 : _GEN_21380; // @[rob.scala 147:39]
  wire  _GEN_25733 = io_i_ex_res_packs_1_valid ? _GEN_23557 : _GEN_21381; // @[rob.scala 147:39]
  wire  _GEN_25734 = io_i_ex_res_packs_1_valid ? _GEN_23558 : _GEN_21382; // @[rob.scala 147:39]
  wire  _GEN_25735 = io_i_ex_res_packs_1_valid ? _GEN_23559 : _GEN_21383; // @[rob.scala 147:39]
  wire  _GEN_25736 = io_i_ex_res_packs_1_valid ? _GEN_23560 : _GEN_21384; // @[rob.scala 147:39]
  wire  _GEN_25737 = io_i_ex_res_packs_1_valid ? _GEN_23561 : _GEN_21385; // @[rob.scala 147:39]
  wire  _GEN_25738 = io_i_ex_res_packs_1_valid ? _GEN_23562 : _GEN_21386; // @[rob.scala 147:39]
  wire  _GEN_25739 = io_i_ex_res_packs_1_valid ? _GEN_23563 : _GEN_21387; // @[rob.scala 147:39]
  wire  _GEN_25740 = io_i_ex_res_packs_1_valid ? _GEN_23564 : _GEN_21388; // @[rob.scala 147:39]
  wire  _GEN_25741 = io_i_ex_res_packs_1_valid ? _GEN_23565 : _GEN_21389; // @[rob.scala 147:39]
  wire  _GEN_25742 = io_i_ex_res_packs_1_valid ? _GEN_23566 : _GEN_21390; // @[rob.scala 147:39]
  wire  _GEN_25743 = io_i_ex_res_packs_1_valid ? _GEN_23567 : _GEN_21391; // @[rob.scala 147:39]
  wire  _GEN_25744 = io_i_ex_res_packs_1_valid ? _GEN_23568 : _GEN_21392; // @[rob.scala 147:39]
  wire  _GEN_25745 = io_i_ex_res_packs_1_valid ? _GEN_23569 : _GEN_21393; // @[rob.scala 147:39]
  wire  _GEN_25746 = io_i_ex_res_packs_1_valid ? _GEN_23570 : _GEN_21394; // @[rob.scala 147:39]
  wire  _GEN_25747 = io_i_ex_res_packs_1_valid ? _GEN_23571 : _GEN_21395; // @[rob.scala 147:39]
  wire  _GEN_25748 = io_i_ex_res_packs_1_valid ? _GEN_23572 : _GEN_21396; // @[rob.scala 147:39]
  wire  _GEN_25749 = io_i_ex_res_packs_1_valid ? _GEN_23573 : _GEN_21397; // @[rob.scala 147:39]
  wire  _GEN_25750 = io_i_ex_res_packs_1_valid ? _GEN_23574 : _GEN_21398; // @[rob.scala 147:39]
  wire  _GEN_25751 = io_i_ex_res_packs_1_valid ? _GEN_23575 : _GEN_21399; // @[rob.scala 147:39]
  wire  _GEN_25752 = io_i_ex_res_packs_1_valid ? _GEN_23576 : _GEN_21400; // @[rob.scala 147:39]
  wire  _GEN_25753 = io_i_ex_res_packs_1_valid ? _GEN_23577 : _GEN_21401; // @[rob.scala 147:39]
  wire  _GEN_25754 = io_i_ex_res_packs_1_valid ? _GEN_23578 : _GEN_21402; // @[rob.scala 147:39]
  wire  _GEN_25755 = io_i_ex_res_packs_1_valid ? _GEN_23579 : _GEN_21403; // @[rob.scala 147:39]
  wire  _GEN_25756 = io_i_ex_res_packs_1_valid ? _GEN_23580 : _GEN_21404; // @[rob.scala 147:39]
  wire  _GEN_25757 = io_i_ex_res_packs_1_valid ? _GEN_23581 : _GEN_21405; // @[rob.scala 147:39]
  wire  _GEN_25758 = io_i_ex_res_packs_1_valid ? _GEN_23582 : _GEN_21406; // @[rob.scala 147:39]
  wire  _GEN_25759 = io_i_ex_res_packs_1_valid ? _GEN_23583 : _GEN_21407; // @[rob.scala 147:39]
  wire  _GEN_25760 = io_i_ex_res_packs_1_valid ? _GEN_23584 : _GEN_21408; // @[rob.scala 147:39]
  wire  _GEN_25761 = io_i_ex_res_packs_1_valid ? _GEN_23585 : _GEN_21409; // @[rob.scala 147:39]
  wire  _GEN_25762 = io_i_ex_res_packs_1_valid ? _GEN_23586 : _GEN_21410; // @[rob.scala 147:39]
  wire  _GEN_25763 = io_i_ex_res_packs_1_valid ? _GEN_23587 : _GEN_21411; // @[rob.scala 147:39]
  wire  _GEN_25764 = io_i_ex_res_packs_1_valid ? _GEN_23588 : _GEN_21412; // @[rob.scala 147:39]
  wire  _GEN_25765 = io_i_ex_res_packs_1_valid ? _GEN_23589 : _GEN_21413; // @[rob.scala 147:39]
  wire  _GEN_25766 = io_i_ex_res_packs_1_valid ? _GEN_23590 : _GEN_21414; // @[rob.scala 147:39]
  wire  _GEN_25767 = io_i_ex_res_packs_1_valid ? _GEN_23591 : _GEN_21415; // @[rob.scala 147:39]
  wire  _GEN_25768 = io_i_ex_res_packs_1_valid ? _GEN_23592 : _GEN_21416; // @[rob.scala 147:39]
  wire  _GEN_25769 = io_i_ex_res_packs_1_valid ? _GEN_23593 : _GEN_21417; // @[rob.scala 147:39]
  wire  _GEN_25770 = io_i_ex_res_packs_1_valid ? _GEN_23594 : _GEN_21418; // @[rob.scala 147:39]
  wire  _GEN_25771 = io_i_ex_res_packs_1_valid ? _GEN_23595 : _GEN_21419; // @[rob.scala 147:39]
  wire  _GEN_25772 = io_i_ex_res_packs_1_valid ? _GEN_23596 : _GEN_21420; // @[rob.scala 147:39]
  wire  _GEN_25773 = io_i_ex_res_packs_1_valid ? _GEN_23597 : _GEN_21421; // @[rob.scala 147:39]
  wire  _GEN_25774 = io_i_ex_res_packs_1_valid ? _GEN_23598 : _GEN_21422; // @[rob.scala 147:39]
  wire  _GEN_25775 = io_i_ex_res_packs_1_valid ? _GEN_23599 : _GEN_21423; // @[rob.scala 147:39]
  wire  _GEN_25776 = io_i_ex_res_packs_1_valid ? _GEN_23600 : _GEN_21424; // @[rob.scala 147:39]
  wire  _GEN_25777 = io_i_ex_res_packs_1_valid ? _GEN_23601 : _GEN_21425; // @[rob.scala 147:39]
  wire  _GEN_25778 = io_i_ex_res_packs_1_valid ? _GEN_23602 : _GEN_21426; // @[rob.scala 147:39]
  wire  _GEN_25779 = io_i_ex_res_packs_1_valid ? _GEN_23603 : _GEN_21427; // @[rob.scala 147:39]
  wire  _GEN_25780 = io_i_ex_res_packs_1_valid ? _GEN_23604 : _GEN_21428; // @[rob.scala 147:39]
  wire  _GEN_25781 = io_i_ex_res_packs_1_valid ? _GEN_23605 : _GEN_21429; // @[rob.scala 147:39]
  wire  _GEN_25782 = io_i_ex_res_packs_1_valid ? _GEN_23606 : _GEN_21430; // @[rob.scala 147:39]
  wire  _GEN_25783 = io_i_ex_res_packs_1_valid ? _GEN_23607 : _GEN_21431; // @[rob.scala 147:39]
  wire  _GEN_25784 = io_i_ex_res_packs_1_valid ? _GEN_23608 : _GEN_21432; // @[rob.scala 147:39]
  wire  _GEN_25785 = io_i_ex_res_packs_1_valid ? _GEN_23609 : _GEN_21433; // @[rob.scala 147:39]
  wire  _GEN_25786 = io_i_ex_res_packs_1_valid ? _GEN_23610 : _GEN_21434; // @[rob.scala 147:39]
  wire  _GEN_25787 = io_i_ex_res_packs_1_valid ? _GEN_23611 : _GEN_21435; // @[rob.scala 147:39]
  wire  _GEN_25788 = io_i_ex_res_packs_1_valid ? _GEN_23612 : _GEN_21436; // @[rob.scala 147:39]
  wire  _GEN_25789 = io_i_ex_res_packs_1_valid ? _GEN_23613 : _GEN_21437; // @[rob.scala 147:39]
  wire  _GEN_25790 = io_i_ex_res_packs_1_valid ? _GEN_23614 : _GEN_21438; // @[rob.scala 147:39]
  wire  _GEN_25791 = io_i_ex_res_packs_1_valid ? _GEN_23615 : _GEN_21439; // @[rob.scala 147:39]
  wire  _GEN_25792 = io_i_ex_res_packs_1_valid ? _GEN_23616 : _GEN_21440; // @[rob.scala 147:39]
  wire  _GEN_25793 = io_i_ex_res_packs_1_valid ? _GEN_23617 : _GEN_21441; // @[rob.scala 147:39]
  wire [31:0] _GEN_25858 = io_i_ex_res_packs_1_valid ? _GEN_23682 : _GEN_21506; // @[rob.scala 147:39]
  wire [31:0] _GEN_25859 = io_i_ex_res_packs_1_valid ? _GEN_23683 : _GEN_21507; // @[rob.scala 147:39]
  wire [31:0] _GEN_25860 = io_i_ex_res_packs_1_valid ? _GEN_23684 : _GEN_21508; // @[rob.scala 147:39]
  wire [31:0] _GEN_25861 = io_i_ex_res_packs_1_valid ? _GEN_23685 : _GEN_21509; // @[rob.scala 147:39]
  wire [31:0] _GEN_25862 = io_i_ex_res_packs_1_valid ? _GEN_23686 : _GEN_21510; // @[rob.scala 147:39]
  wire [31:0] _GEN_25863 = io_i_ex_res_packs_1_valid ? _GEN_23687 : _GEN_21511; // @[rob.scala 147:39]
  wire [31:0] _GEN_25864 = io_i_ex_res_packs_1_valid ? _GEN_23688 : _GEN_21512; // @[rob.scala 147:39]
  wire [31:0] _GEN_25865 = io_i_ex_res_packs_1_valid ? _GEN_23689 : _GEN_21513; // @[rob.scala 147:39]
  wire [31:0] _GEN_25866 = io_i_ex_res_packs_1_valid ? _GEN_23690 : _GEN_21514; // @[rob.scala 147:39]
  wire [31:0] _GEN_25867 = io_i_ex_res_packs_1_valid ? _GEN_23691 : _GEN_21515; // @[rob.scala 147:39]
  wire [31:0] _GEN_25868 = io_i_ex_res_packs_1_valid ? _GEN_23692 : _GEN_21516; // @[rob.scala 147:39]
  wire [31:0] _GEN_25869 = io_i_ex_res_packs_1_valid ? _GEN_23693 : _GEN_21517; // @[rob.scala 147:39]
  wire [31:0] _GEN_25870 = io_i_ex_res_packs_1_valid ? _GEN_23694 : _GEN_21518; // @[rob.scala 147:39]
  wire [31:0] _GEN_25871 = io_i_ex_res_packs_1_valid ? _GEN_23695 : _GEN_21519; // @[rob.scala 147:39]
  wire [31:0] _GEN_25872 = io_i_ex_res_packs_1_valid ? _GEN_23696 : _GEN_21520; // @[rob.scala 147:39]
  wire [31:0] _GEN_25873 = io_i_ex_res_packs_1_valid ? _GEN_23697 : _GEN_21521; // @[rob.scala 147:39]
  wire [31:0] _GEN_25874 = io_i_ex_res_packs_1_valid ? _GEN_23698 : _GEN_21522; // @[rob.scala 147:39]
  wire [31:0] _GEN_25875 = io_i_ex_res_packs_1_valid ? _GEN_23699 : _GEN_21523; // @[rob.scala 147:39]
  wire [31:0] _GEN_25876 = io_i_ex_res_packs_1_valid ? _GEN_23700 : _GEN_21524; // @[rob.scala 147:39]
  wire [31:0] _GEN_25877 = io_i_ex_res_packs_1_valid ? _GEN_23701 : _GEN_21525; // @[rob.scala 147:39]
  wire [31:0] _GEN_25878 = io_i_ex_res_packs_1_valid ? _GEN_23702 : _GEN_21526; // @[rob.scala 147:39]
  wire [31:0] _GEN_25879 = io_i_ex_res_packs_1_valid ? _GEN_23703 : _GEN_21527; // @[rob.scala 147:39]
  wire [31:0] _GEN_25880 = io_i_ex_res_packs_1_valid ? _GEN_23704 : _GEN_21528; // @[rob.scala 147:39]
  wire [31:0] _GEN_25881 = io_i_ex_res_packs_1_valid ? _GEN_23705 : _GEN_21529; // @[rob.scala 147:39]
  wire [31:0] _GEN_25882 = io_i_ex_res_packs_1_valid ? _GEN_23706 : _GEN_21530; // @[rob.scala 147:39]
  wire [31:0] _GEN_25883 = io_i_ex_res_packs_1_valid ? _GEN_23707 : _GEN_21531; // @[rob.scala 147:39]
  wire [31:0] _GEN_25884 = io_i_ex_res_packs_1_valid ? _GEN_23708 : _GEN_21532; // @[rob.scala 147:39]
  wire [31:0] _GEN_25885 = io_i_ex_res_packs_1_valid ? _GEN_23709 : _GEN_21533; // @[rob.scala 147:39]
  wire [31:0] _GEN_25886 = io_i_ex_res_packs_1_valid ? _GEN_23710 : _GEN_21534; // @[rob.scala 147:39]
  wire [31:0] _GEN_25887 = io_i_ex_res_packs_1_valid ? _GEN_23711 : _GEN_21535; // @[rob.scala 147:39]
  wire [31:0] _GEN_25888 = io_i_ex_res_packs_1_valid ? _GEN_23712 : _GEN_21536; // @[rob.scala 147:39]
  wire [31:0] _GEN_25889 = io_i_ex_res_packs_1_valid ? _GEN_23713 : _GEN_21537; // @[rob.scala 147:39]
  wire [31:0] _GEN_25890 = io_i_ex_res_packs_1_valid ? _GEN_23714 : _GEN_21538; // @[rob.scala 147:39]
  wire [31:0] _GEN_25891 = io_i_ex_res_packs_1_valid ? _GEN_23715 : _GEN_21539; // @[rob.scala 147:39]
  wire [31:0] _GEN_25892 = io_i_ex_res_packs_1_valid ? _GEN_23716 : _GEN_21540; // @[rob.scala 147:39]
  wire [31:0] _GEN_25893 = io_i_ex_res_packs_1_valid ? _GEN_23717 : _GEN_21541; // @[rob.scala 147:39]
  wire [31:0] _GEN_25894 = io_i_ex_res_packs_1_valid ? _GEN_23718 : _GEN_21542; // @[rob.scala 147:39]
  wire [31:0] _GEN_25895 = io_i_ex_res_packs_1_valid ? _GEN_23719 : _GEN_21543; // @[rob.scala 147:39]
  wire [31:0] _GEN_25896 = io_i_ex_res_packs_1_valid ? _GEN_23720 : _GEN_21544; // @[rob.scala 147:39]
  wire [31:0] _GEN_25897 = io_i_ex_res_packs_1_valid ? _GEN_23721 : _GEN_21545; // @[rob.scala 147:39]
  wire [31:0] _GEN_25898 = io_i_ex_res_packs_1_valid ? _GEN_23722 : _GEN_21546; // @[rob.scala 147:39]
  wire [31:0] _GEN_25899 = io_i_ex_res_packs_1_valid ? _GEN_23723 : _GEN_21547; // @[rob.scala 147:39]
  wire [31:0] _GEN_25900 = io_i_ex_res_packs_1_valid ? _GEN_23724 : _GEN_21548; // @[rob.scala 147:39]
  wire [31:0] _GEN_25901 = io_i_ex_res_packs_1_valid ? _GEN_23725 : _GEN_21549; // @[rob.scala 147:39]
  wire [31:0] _GEN_25902 = io_i_ex_res_packs_1_valid ? _GEN_23726 : _GEN_21550; // @[rob.scala 147:39]
  wire [31:0] _GEN_25903 = io_i_ex_res_packs_1_valid ? _GEN_23727 : _GEN_21551; // @[rob.scala 147:39]
  wire [31:0] _GEN_25904 = io_i_ex_res_packs_1_valid ? _GEN_23728 : _GEN_21552; // @[rob.scala 147:39]
  wire [31:0] _GEN_25905 = io_i_ex_res_packs_1_valid ? _GEN_23729 : _GEN_21553; // @[rob.scala 147:39]
  wire [31:0] _GEN_25906 = io_i_ex_res_packs_1_valid ? _GEN_23730 : _GEN_21554; // @[rob.scala 147:39]
  wire [31:0] _GEN_25907 = io_i_ex_res_packs_1_valid ? _GEN_23731 : _GEN_21555; // @[rob.scala 147:39]
  wire [31:0] _GEN_25908 = io_i_ex_res_packs_1_valid ? _GEN_23732 : _GEN_21556; // @[rob.scala 147:39]
  wire [31:0] _GEN_25909 = io_i_ex_res_packs_1_valid ? _GEN_23733 : _GEN_21557; // @[rob.scala 147:39]
  wire [31:0] _GEN_25910 = io_i_ex_res_packs_1_valid ? _GEN_23734 : _GEN_21558; // @[rob.scala 147:39]
  wire [31:0] _GEN_25911 = io_i_ex_res_packs_1_valid ? _GEN_23735 : _GEN_21559; // @[rob.scala 147:39]
  wire [31:0] _GEN_25912 = io_i_ex_res_packs_1_valid ? _GEN_23736 : _GEN_21560; // @[rob.scala 147:39]
  wire [31:0] _GEN_25913 = io_i_ex_res_packs_1_valid ? _GEN_23737 : _GEN_21561; // @[rob.scala 147:39]
  wire [31:0] _GEN_25914 = io_i_ex_res_packs_1_valid ? _GEN_23738 : _GEN_21562; // @[rob.scala 147:39]
  wire [31:0] _GEN_25915 = io_i_ex_res_packs_1_valid ? _GEN_23739 : _GEN_21563; // @[rob.scala 147:39]
  wire [31:0] _GEN_25916 = io_i_ex_res_packs_1_valid ? _GEN_23740 : _GEN_21564; // @[rob.scala 147:39]
  wire [31:0] _GEN_25917 = io_i_ex_res_packs_1_valid ? _GEN_23741 : _GEN_21565; // @[rob.scala 147:39]
  wire [31:0] _GEN_25918 = io_i_ex_res_packs_1_valid ? _GEN_23742 : _GEN_21566; // @[rob.scala 147:39]
  wire [31:0] _GEN_25919 = io_i_ex_res_packs_1_valid ? _GEN_23743 : _GEN_21567; // @[rob.scala 147:39]
  wire [31:0] _GEN_25920 = io_i_ex_res_packs_1_valid ? _GEN_23744 : _GEN_21568; // @[rob.scala 147:39]
  wire [31:0] _GEN_25921 = io_i_ex_res_packs_1_valid ? _GEN_23745 : _GEN_21569; // @[rob.scala 147:39]
  wire [31:0] _GEN_25922 = io_i_ex_res_packs_1_valid ? _GEN_23746 : _GEN_21570; // @[rob.scala 147:39]
  wire [31:0] _GEN_25923 = io_i_ex_res_packs_1_valid ? _GEN_23747 : _GEN_21571; // @[rob.scala 147:39]
  wire [31:0] _GEN_25924 = io_i_ex_res_packs_1_valid ? _GEN_23748 : _GEN_21572; // @[rob.scala 147:39]
  wire [31:0] _GEN_25925 = io_i_ex_res_packs_1_valid ? _GEN_23749 : _GEN_21573; // @[rob.scala 147:39]
  wire [31:0] _GEN_25926 = io_i_ex_res_packs_1_valid ? _GEN_23750 : _GEN_21574; // @[rob.scala 147:39]
  wire [31:0] _GEN_25927 = io_i_ex_res_packs_1_valid ? _GEN_23751 : _GEN_21575; // @[rob.scala 147:39]
  wire [31:0] _GEN_25928 = io_i_ex_res_packs_1_valid ? _GEN_23752 : _GEN_21576; // @[rob.scala 147:39]
  wire [31:0] _GEN_25929 = io_i_ex_res_packs_1_valid ? _GEN_23753 : _GEN_21577; // @[rob.scala 147:39]
  wire [31:0] _GEN_25930 = io_i_ex_res_packs_1_valid ? _GEN_23754 : _GEN_21578; // @[rob.scala 147:39]
  wire [31:0] _GEN_25931 = io_i_ex_res_packs_1_valid ? _GEN_23755 : _GEN_21579; // @[rob.scala 147:39]
  wire [31:0] _GEN_25932 = io_i_ex_res_packs_1_valid ? _GEN_23756 : _GEN_21580; // @[rob.scala 147:39]
  wire [31:0] _GEN_25933 = io_i_ex_res_packs_1_valid ? _GEN_23757 : _GEN_21581; // @[rob.scala 147:39]
  wire [31:0] _GEN_25934 = io_i_ex_res_packs_1_valid ? _GEN_23758 : _GEN_21582; // @[rob.scala 147:39]
  wire [31:0] _GEN_25935 = io_i_ex_res_packs_1_valid ? _GEN_23759 : _GEN_21583; // @[rob.scala 147:39]
  wire [31:0] _GEN_25936 = io_i_ex_res_packs_1_valid ? _GEN_23760 : _GEN_21584; // @[rob.scala 147:39]
  wire [31:0] _GEN_25937 = io_i_ex_res_packs_1_valid ? _GEN_23761 : _GEN_21585; // @[rob.scala 147:39]
  wire [31:0] _GEN_25938 = io_i_ex_res_packs_1_valid ? _GEN_23762 : _GEN_21586; // @[rob.scala 147:39]
  wire [31:0] _GEN_25939 = io_i_ex_res_packs_1_valid ? _GEN_23763 : _GEN_21587; // @[rob.scala 147:39]
  wire [31:0] _GEN_25940 = io_i_ex_res_packs_1_valid ? _GEN_23764 : _GEN_21588; // @[rob.scala 147:39]
  wire [31:0] _GEN_25941 = io_i_ex_res_packs_1_valid ? _GEN_23765 : _GEN_21589; // @[rob.scala 147:39]
  wire [31:0] _GEN_25942 = io_i_ex_res_packs_1_valid ? _GEN_23766 : _GEN_21590; // @[rob.scala 147:39]
  wire [31:0] _GEN_25943 = io_i_ex_res_packs_1_valid ? _GEN_23767 : _GEN_21591; // @[rob.scala 147:39]
  wire [31:0] _GEN_25944 = io_i_ex_res_packs_1_valid ? _GEN_23768 : _GEN_21592; // @[rob.scala 147:39]
  wire [31:0] _GEN_25945 = io_i_ex_res_packs_1_valid ? _GEN_23769 : _GEN_21593; // @[rob.scala 147:39]
  wire [31:0] _GEN_25946 = io_i_ex_res_packs_1_valid ? _GEN_23770 : _GEN_21594; // @[rob.scala 147:39]
  wire [31:0] _GEN_25947 = io_i_ex_res_packs_1_valid ? _GEN_23771 : _GEN_21595; // @[rob.scala 147:39]
  wire [31:0] _GEN_25948 = io_i_ex_res_packs_1_valid ? _GEN_23772 : _GEN_21596; // @[rob.scala 147:39]
  wire [31:0] _GEN_25949 = io_i_ex_res_packs_1_valid ? _GEN_23773 : _GEN_21597; // @[rob.scala 147:39]
  wire [31:0] _GEN_25950 = io_i_ex_res_packs_1_valid ? _GEN_23774 : _GEN_21598; // @[rob.scala 147:39]
  wire [31:0] _GEN_25951 = io_i_ex_res_packs_1_valid ? _GEN_23775 : _GEN_21599; // @[rob.scala 147:39]
  wire [31:0] _GEN_25952 = io_i_ex_res_packs_1_valid ? _GEN_23776 : _GEN_21600; // @[rob.scala 147:39]
  wire [31:0] _GEN_25953 = io_i_ex_res_packs_1_valid ? _GEN_23777 : _GEN_21601; // @[rob.scala 147:39]
  wire [31:0] _GEN_25954 = io_i_ex_res_packs_1_valid ? _GEN_23778 : _GEN_21602; // @[rob.scala 147:39]
  wire [31:0] _GEN_25955 = io_i_ex_res_packs_1_valid ? _GEN_23779 : _GEN_21603; // @[rob.scala 147:39]
  wire [31:0] _GEN_25956 = io_i_ex_res_packs_1_valid ? _GEN_23780 : _GEN_21604; // @[rob.scala 147:39]
  wire [31:0] _GEN_25957 = io_i_ex_res_packs_1_valid ? _GEN_23781 : _GEN_21605; // @[rob.scala 147:39]
  wire [31:0] _GEN_25958 = io_i_ex_res_packs_1_valid ? _GEN_23782 : _GEN_21606; // @[rob.scala 147:39]
  wire [31:0] _GEN_25959 = io_i_ex_res_packs_1_valid ? _GEN_23783 : _GEN_21607; // @[rob.scala 147:39]
  wire [31:0] _GEN_25960 = io_i_ex_res_packs_1_valid ? _GEN_23784 : _GEN_21608; // @[rob.scala 147:39]
  wire [31:0] _GEN_25961 = io_i_ex_res_packs_1_valid ? _GEN_23785 : _GEN_21609; // @[rob.scala 147:39]
  wire [31:0] _GEN_25962 = io_i_ex_res_packs_1_valid ? _GEN_23786 : _GEN_21610; // @[rob.scala 147:39]
  wire [31:0] _GEN_25963 = io_i_ex_res_packs_1_valid ? _GEN_23787 : _GEN_21611; // @[rob.scala 147:39]
  wire [31:0] _GEN_25964 = io_i_ex_res_packs_1_valid ? _GEN_23788 : _GEN_21612; // @[rob.scala 147:39]
  wire [31:0] _GEN_25965 = io_i_ex_res_packs_1_valid ? _GEN_23789 : _GEN_21613; // @[rob.scala 147:39]
  wire [31:0] _GEN_25966 = io_i_ex_res_packs_1_valid ? _GEN_23790 : _GEN_21614; // @[rob.scala 147:39]
  wire [31:0] _GEN_25967 = io_i_ex_res_packs_1_valid ? _GEN_23791 : _GEN_21615; // @[rob.scala 147:39]
  wire [31:0] _GEN_25968 = io_i_ex_res_packs_1_valid ? _GEN_23792 : _GEN_21616; // @[rob.scala 147:39]
  wire [31:0] _GEN_25969 = io_i_ex_res_packs_1_valid ? _GEN_23793 : _GEN_21617; // @[rob.scala 147:39]
  wire [31:0] _GEN_25970 = io_i_ex_res_packs_1_valid ? _GEN_23794 : _GEN_21618; // @[rob.scala 147:39]
  wire [31:0] _GEN_25971 = io_i_ex_res_packs_1_valid ? _GEN_23795 : _GEN_21619; // @[rob.scala 147:39]
  wire [31:0] _GEN_25972 = io_i_ex_res_packs_1_valid ? _GEN_23796 : _GEN_21620; // @[rob.scala 147:39]
  wire [31:0] _GEN_25973 = io_i_ex_res_packs_1_valid ? _GEN_23797 : _GEN_21621; // @[rob.scala 147:39]
  wire [31:0] _GEN_25974 = io_i_ex_res_packs_1_valid ? _GEN_23798 : _GEN_21622; // @[rob.scala 147:39]
  wire [31:0] _GEN_25975 = io_i_ex_res_packs_1_valid ? _GEN_23799 : _GEN_21623; // @[rob.scala 147:39]
  wire [31:0] _GEN_25976 = io_i_ex_res_packs_1_valid ? _GEN_23800 : _GEN_21624; // @[rob.scala 147:39]
  wire [31:0] _GEN_25977 = io_i_ex_res_packs_1_valid ? _GEN_23801 : _GEN_21625; // @[rob.scala 147:39]
  wire [31:0] _GEN_25978 = io_i_ex_res_packs_1_valid ? _GEN_23802 : _GEN_21626; // @[rob.scala 147:39]
  wire [31:0] _GEN_25979 = io_i_ex_res_packs_1_valid ? _GEN_23803 : _GEN_21627; // @[rob.scala 147:39]
  wire [31:0] _GEN_25980 = io_i_ex_res_packs_1_valid ? _GEN_23804 : _GEN_21628; // @[rob.scala 147:39]
  wire [31:0] _GEN_25981 = io_i_ex_res_packs_1_valid ? _GEN_23805 : _GEN_21629; // @[rob.scala 147:39]
  wire [31:0] _GEN_25982 = io_i_ex_res_packs_1_valid ? _GEN_23806 : _GEN_21630; // @[rob.scala 147:39]
  wire [31:0] _GEN_25983 = io_i_ex_res_packs_1_valid ? _GEN_23807 : _GEN_21631; // @[rob.scala 147:39]
  wire [31:0] _GEN_25984 = io_i_ex_res_packs_1_valid ? _GEN_23808 : _GEN_21632; // @[rob.scala 147:39]
  wire [31:0] _GEN_25985 = io_i_ex_res_packs_1_valid ? _GEN_23809 : _GEN_21633; // @[rob.scala 147:39]
  wire [6:0] _GEN_25986 = io_i_ex_res_packs_1_valid ? _GEN_23810 : _GEN_21634; // @[rob.scala 147:39]
  wire [6:0] _GEN_25987 = io_i_ex_res_packs_1_valid ? _GEN_23811 : _GEN_21635; // @[rob.scala 147:39]
  wire [6:0] _GEN_25988 = io_i_ex_res_packs_1_valid ? _GEN_23812 : _GEN_21636; // @[rob.scala 147:39]
  wire [6:0] _GEN_25989 = io_i_ex_res_packs_1_valid ? _GEN_23813 : _GEN_21637; // @[rob.scala 147:39]
  wire [6:0] _GEN_25990 = io_i_ex_res_packs_1_valid ? _GEN_23814 : _GEN_21638; // @[rob.scala 147:39]
  wire [6:0] _GEN_25991 = io_i_ex_res_packs_1_valid ? _GEN_23815 : _GEN_21639; // @[rob.scala 147:39]
  wire [6:0] _GEN_25992 = io_i_ex_res_packs_1_valid ? _GEN_23816 : _GEN_21640; // @[rob.scala 147:39]
  wire [6:0] _GEN_25993 = io_i_ex_res_packs_1_valid ? _GEN_23817 : _GEN_21641; // @[rob.scala 147:39]
  wire [6:0] _GEN_25994 = io_i_ex_res_packs_1_valid ? _GEN_23818 : _GEN_21642; // @[rob.scala 147:39]
  wire [6:0] _GEN_25995 = io_i_ex_res_packs_1_valid ? _GEN_23819 : _GEN_21643; // @[rob.scala 147:39]
  wire [6:0] _GEN_25996 = io_i_ex_res_packs_1_valid ? _GEN_23820 : _GEN_21644; // @[rob.scala 147:39]
  wire [6:0] _GEN_25997 = io_i_ex_res_packs_1_valid ? _GEN_23821 : _GEN_21645; // @[rob.scala 147:39]
  wire [6:0] _GEN_25998 = io_i_ex_res_packs_1_valid ? _GEN_23822 : _GEN_21646; // @[rob.scala 147:39]
  wire [6:0] _GEN_25999 = io_i_ex_res_packs_1_valid ? _GEN_23823 : _GEN_21647; // @[rob.scala 147:39]
  wire [6:0] _GEN_26000 = io_i_ex_res_packs_1_valid ? _GEN_23824 : _GEN_21648; // @[rob.scala 147:39]
  wire [6:0] _GEN_26001 = io_i_ex_res_packs_1_valid ? _GEN_23825 : _GEN_21649; // @[rob.scala 147:39]
  wire [6:0] _GEN_26002 = io_i_ex_res_packs_1_valid ? _GEN_23826 : _GEN_21650; // @[rob.scala 147:39]
  wire [6:0] _GEN_26003 = io_i_ex_res_packs_1_valid ? _GEN_23827 : _GEN_21651; // @[rob.scala 147:39]
  wire [6:0] _GEN_26004 = io_i_ex_res_packs_1_valid ? _GEN_23828 : _GEN_21652; // @[rob.scala 147:39]
  wire [6:0] _GEN_26005 = io_i_ex_res_packs_1_valid ? _GEN_23829 : _GEN_21653; // @[rob.scala 147:39]
  wire [6:0] _GEN_26006 = io_i_ex_res_packs_1_valid ? _GEN_23830 : _GEN_21654; // @[rob.scala 147:39]
  wire [6:0] _GEN_26007 = io_i_ex_res_packs_1_valid ? _GEN_23831 : _GEN_21655; // @[rob.scala 147:39]
  wire [6:0] _GEN_26008 = io_i_ex_res_packs_1_valid ? _GEN_23832 : _GEN_21656; // @[rob.scala 147:39]
  wire [6:0] _GEN_26009 = io_i_ex_res_packs_1_valid ? _GEN_23833 : _GEN_21657; // @[rob.scala 147:39]
  wire [6:0] _GEN_26010 = io_i_ex_res_packs_1_valid ? _GEN_23834 : _GEN_21658; // @[rob.scala 147:39]
  wire [6:0] _GEN_26011 = io_i_ex_res_packs_1_valid ? _GEN_23835 : _GEN_21659; // @[rob.scala 147:39]
  wire [6:0] _GEN_26012 = io_i_ex_res_packs_1_valid ? _GEN_23836 : _GEN_21660; // @[rob.scala 147:39]
  wire [6:0] _GEN_26013 = io_i_ex_res_packs_1_valid ? _GEN_23837 : _GEN_21661; // @[rob.scala 147:39]
  wire [6:0] _GEN_26014 = io_i_ex_res_packs_1_valid ? _GEN_23838 : _GEN_21662; // @[rob.scala 147:39]
  wire [6:0] _GEN_26015 = io_i_ex_res_packs_1_valid ? _GEN_23839 : _GEN_21663; // @[rob.scala 147:39]
  wire [6:0] _GEN_26016 = io_i_ex_res_packs_1_valid ? _GEN_23840 : _GEN_21664; // @[rob.scala 147:39]
  wire [6:0] _GEN_26017 = io_i_ex_res_packs_1_valid ? _GEN_23841 : _GEN_21665; // @[rob.scala 147:39]
  wire [6:0] _GEN_26018 = io_i_ex_res_packs_1_valid ? _GEN_23842 : _GEN_21666; // @[rob.scala 147:39]
  wire [6:0] _GEN_26019 = io_i_ex_res_packs_1_valid ? _GEN_23843 : _GEN_21667; // @[rob.scala 147:39]
  wire [6:0] _GEN_26020 = io_i_ex_res_packs_1_valid ? _GEN_23844 : _GEN_21668; // @[rob.scala 147:39]
  wire [6:0] _GEN_26021 = io_i_ex_res_packs_1_valid ? _GEN_23845 : _GEN_21669; // @[rob.scala 147:39]
  wire [6:0] _GEN_26022 = io_i_ex_res_packs_1_valid ? _GEN_23846 : _GEN_21670; // @[rob.scala 147:39]
  wire [6:0] _GEN_26023 = io_i_ex_res_packs_1_valid ? _GEN_23847 : _GEN_21671; // @[rob.scala 147:39]
  wire [6:0] _GEN_26024 = io_i_ex_res_packs_1_valid ? _GEN_23848 : _GEN_21672; // @[rob.scala 147:39]
  wire [6:0] _GEN_26025 = io_i_ex_res_packs_1_valid ? _GEN_23849 : _GEN_21673; // @[rob.scala 147:39]
  wire [6:0] _GEN_26026 = io_i_ex_res_packs_1_valid ? _GEN_23850 : _GEN_21674; // @[rob.scala 147:39]
  wire [6:0] _GEN_26027 = io_i_ex_res_packs_1_valid ? _GEN_23851 : _GEN_21675; // @[rob.scala 147:39]
  wire [6:0] _GEN_26028 = io_i_ex_res_packs_1_valid ? _GEN_23852 : _GEN_21676; // @[rob.scala 147:39]
  wire [6:0] _GEN_26029 = io_i_ex_res_packs_1_valid ? _GEN_23853 : _GEN_21677; // @[rob.scala 147:39]
  wire [6:0] _GEN_26030 = io_i_ex_res_packs_1_valid ? _GEN_23854 : _GEN_21678; // @[rob.scala 147:39]
  wire [6:0] _GEN_26031 = io_i_ex_res_packs_1_valid ? _GEN_23855 : _GEN_21679; // @[rob.scala 147:39]
  wire [6:0] _GEN_26032 = io_i_ex_res_packs_1_valid ? _GEN_23856 : _GEN_21680; // @[rob.scala 147:39]
  wire [6:0] _GEN_26033 = io_i_ex_res_packs_1_valid ? _GEN_23857 : _GEN_21681; // @[rob.scala 147:39]
  wire [6:0] _GEN_26034 = io_i_ex_res_packs_1_valid ? _GEN_23858 : _GEN_21682; // @[rob.scala 147:39]
  wire [6:0] _GEN_26035 = io_i_ex_res_packs_1_valid ? _GEN_23859 : _GEN_21683; // @[rob.scala 147:39]
  wire [6:0] _GEN_26036 = io_i_ex_res_packs_1_valid ? _GEN_23860 : _GEN_21684; // @[rob.scala 147:39]
  wire [6:0] _GEN_26037 = io_i_ex_res_packs_1_valid ? _GEN_23861 : _GEN_21685; // @[rob.scala 147:39]
  wire [6:0] _GEN_26038 = io_i_ex_res_packs_1_valid ? _GEN_23862 : _GEN_21686; // @[rob.scala 147:39]
  wire [6:0] _GEN_26039 = io_i_ex_res_packs_1_valid ? _GEN_23863 : _GEN_21687; // @[rob.scala 147:39]
  wire [6:0] _GEN_26040 = io_i_ex_res_packs_1_valid ? _GEN_23864 : _GEN_21688; // @[rob.scala 147:39]
  wire [6:0] _GEN_26041 = io_i_ex_res_packs_1_valid ? _GEN_23865 : _GEN_21689; // @[rob.scala 147:39]
  wire [6:0] _GEN_26042 = io_i_ex_res_packs_1_valid ? _GEN_23866 : _GEN_21690; // @[rob.scala 147:39]
  wire [6:0] _GEN_26043 = io_i_ex_res_packs_1_valid ? _GEN_23867 : _GEN_21691; // @[rob.scala 147:39]
  wire [6:0] _GEN_26044 = io_i_ex_res_packs_1_valid ? _GEN_23868 : _GEN_21692; // @[rob.scala 147:39]
  wire [6:0] _GEN_26045 = io_i_ex_res_packs_1_valid ? _GEN_23869 : _GEN_21693; // @[rob.scala 147:39]
  wire [6:0] _GEN_26046 = io_i_ex_res_packs_1_valid ? _GEN_23870 : _GEN_21694; // @[rob.scala 147:39]
  wire [6:0] _GEN_26047 = io_i_ex_res_packs_1_valid ? _GEN_23871 : _GEN_21695; // @[rob.scala 147:39]
  wire [6:0] _GEN_26048 = io_i_ex_res_packs_1_valid ? _GEN_23872 : _GEN_21696; // @[rob.scala 147:39]
  wire [6:0] _GEN_26049 = io_i_ex_res_packs_1_valid ? _GEN_23873 : _GEN_21697; // @[rob.scala 147:39]
  wire [6:0] _GEN_26370 = io_i_ex_res_packs_1_valid ? _GEN_24194 : _GEN_22018; // @[rob.scala 147:39]
  wire [6:0] _GEN_26371 = io_i_ex_res_packs_1_valid ? _GEN_24195 : _GEN_22019; // @[rob.scala 147:39]
  wire [6:0] _GEN_26372 = io_i_ex_res_packs_1_valid ? _GEN_24196 : _GEN_22020; // @[rob.scala 147:39]
  wire [6:0] _GEN_26373 = io_i_ex_res_packs_1_valid ? _GEN_24197 : _GEN_22021; // @[rob.scala 147:39]
  wire [6:0] _GEN_26374 = io_i_ex_res_packs_1_valid ? _GEN_24198 : _GEN_22022; // @[rob.scala 147:39]
  wire [6:0] _GEN_26375 = io_i_ex_res_packs_1_valid ? _GEN_24199 : _GEN_22023; // @[rob.scala 147:39]
  wire [6:0] _GEN_26376 = io_i_ex_res_packs_1_valid ? _GEN_24200 : _GEN_22024; // @[rob.scala 147:39]
  wire [6:0] _GEN_26377 = io_i_ex_res_packs_1_valid ? _GEN_24201 : _GEN_22025; // @[rob.scala 147:39]
  wire [6:0] _GEN_26378 = io_i_ex_res_packs_1_valid ? _GEN_24202 : _GEN_22026; // @[rob.scala 147:39]
  wire [6:0] _GEN_26379 = io_i_ex_res_packs_1_valid ? _GEN_24203 : _GEN_22027; // @[rob.scala 147:39]
  wire [6:0] _GEN_26380 = io_i_ex_res_packs_1_valid ? _GEN_24204 : _GEN_22028; // @[rob.scala 147:39]
  wire [6:0] _GEN_26381 = io_i_ex_res_packs_1_valid ? _GEN_24205 : _GEN_22029; // @[rob.scala 147:39]
  wire [6:0] _GEN_26382 = io_i_ex_res_packs_1_valid ? _GEN_24206 : _GEN_22030; // @[rob.scala 147:39]
  wire [6:0] _GEN_26383 = io_i_ex_res_packs_1_valid ? _GEN_24207 : _GEN_22031; // @[rob.scala 147:39]
  wire [6:0] _GEN_26384 = io_i_ex_res_packs_1_valid ? _GEN_24208 : _GEN_22032; // @[rob.scala 147:39]
  wire [6:0] _GEN_26385 = io_i_ex_res_packs_1_valid ? _GEN_24209 : _GEN_22033; // @[rob.scala 147:39]
  wire [6:0] _GEN_26386 = io_i_ex_res_packs_1_valid ? _GEN_24210 : _GEN_22034; // @[rob.scala 147:39]
  wire [6:0] _GEN_26387 = io_i_ex_res_packs_1_valid ? _GEN_24211 : _GEN_22035; // @[rob.scala 147:39]
  wire [6:0] _GEN_26388 = io_i_ex_res_packs_1_valid ? _GEN_24212 : _GEN_22036; // @[rob.scala 147:39]
  wire [6:0] _GEN_26389 = io_i_ex_res_packs_1_valid ? _GEN_24213 : _GEN_22037; // @[rob.scala 147:39]
  wire [6:0] _GEN_26390 = io_i_ex_res_packs_1_valid ? _GEN_24214 : _GEN_22038; // @[rob.scala 147:39]
  wire [6:0] _GEN_26391 = io_i_ex_res_packs_1_valid ? _GEN_24215 : _GEN_22039; // @[rob.scala 147:39]
  wire [6:0] _GEN_26392 = io_i_ex_res_packs_1_valid ? _GEN_24216 : _GEN_22040; // @[rob.scala 147:39]
  wire [6:0] _GEN_26393 = io_i_ex_res_packs_1_valid ? _GEN_24217 : _GEN_22041; // @[rob.scala 147:39]
  wire [6:0] _GEN_26394 = io_i_ex_res_packs_1_valid ? _GEN_24218 : _GEN_22042; // @[rob.scala 147:39]
  wire [6:0] _GEN_26395 = io_i_ex_res_packs_1_valid ? _GEN_24219 : _GEN_22043; // @[rob.scala 147:39]
  wire [6:0] _GEN_26396 = io_i_ex_res_packs_1_valid ? _GEN_24220 : _GEN_22044; // @[rob.scala 147:39]
  wire [6:0] _GEN_26397 = io_i_ex_res_packs_1_valid ? _GEN_24221 : _GEN_22045; // @[rob.scala 147:39]
  wire [6:0] _GEN_26398 = io_i_ex_res_packs_1_valid ? _GEN_24222 : _GEN_22046; // @[rob.scala 147:39]
  wire [6:0] _GEN_26399 = io_i_ex_res_packs_1_valid ? _GEN_24223 : _GEN_22047; // @[rob.scala 147:39]
  wire [6:0] _GEN_26400 = io_i_ex_res_packs_1_valid ? _GEN_24224 : _GEN_22048; // @[rob.scala 147:39]
  wire [6:0] _GEN_26401 = io_i_ex_res_packs_1_valid ? _GEN_24225 : _GEN_22049; // @[rob.scala 147:39]
  wire [6:0] _GEN_26402 = io_i_ex_res_packs_1_valid ? _GEN_24226 : _GEN_22050; // @[rob.scala 147:39]
  wire [6:0] _GEN_26403 = io_i_ex_res_packs_1_valid ? _GEN_24227 : _GEN_22051; // @[rob.scala 147:39]
  wire [6:0] _GEN_26404 = io_i_ex_res_packs_1_valid ? _GEN_24228 : _GEN_22052; // @[rob.scala 147:39]
  wire [6:0] _GEN_26405 = io_i_ex_res_packs_1_valid ? _GEN_24229 : _GEN_22053; // @[rob.scala 147:39]
  wire [6:0] _GEN_26406 = io_i_ex_res_packs_1_valid ? _GEN_24230 : _GEN_22054; // @[rob.scala 147:39]
  wire [6:0] _GEN_26407 = io_i_ex_res_packs_1_valid ? _GEN_24231 : _GEN_22055; // @[rob.scala 147:39]
  wire [6:0] _GEN_26408 = io_i_ex_res_packs_1_valid ? _GEN_24232 : _GEN_22056; // @[rob.scala 147:39]
  wire [6:0] _GEN_26409 = io_i_ex_res_packs_1_valid ? _GEN_24233 : _GEN_22057; // @[rob.scala 147:39]
  wire [6:0] _GEN_26410 = io_i_ex_res_packs_1_valid ? _GEN_24234 : _GEN_22058; // @[rob.scala 147:39]
  wire [6:0] _GEN_26411 = io_i_ex_res_packs_1_valid ? _GEN_24235 : _GEN_22059; // @[rob.scala 147:39]
  wire [6:0] _GEN_26412 = io_i_ex_res_packs_1_valid ? _GEN_24236 : _GEN_22060; // @[rob.scala 147:39]
  wire [6:0] _GEN_26413 = io_i_ex_res_packs_1_valid ? _GEN_24237 : _GEN_22061; // @[rob.scala 147:39]
  wire [6:0] _GEN_26414 = io_i_ex_res_packs_1_valid ? _GEN_24238 : _GEN_22062; // @[rob.scala 147:39]
  wire [6:0] _GEN_26415 = io_i_ex_res_packs_1_valid ? _GEN_24239 : _GEN_22063; // @[rob.scala 147:39]
  wire [6:0] _GEN_26416 = io_i_ex_res_packs_1_valid ? _GEN_24240 : _GEN_22064; // @[rob.scala 147:39]
  wire [6:0] _GEN_26417 = io_i_ex_res_packs_1_valid ? _GEN_24241 : _GEN_22065; // @[rob.scala 147:39]
  wire [6:0] _GEN_26418 = io_i_ex_res_packs_1_valid ? _GEN_24242 : _GEN_22066; // @[rob.scala 147:39]
  wire [6:0] _GEN_26419 = io_i_ex_res_packs_1_valid ? _GEN_24243 : _GEN_22067; // @[rob.scala 147:39]
  wire [6:0] _GEN_26420 = io_i_ex_res_packs_1_valid ? _GEN_24244 : _GEN_22068; // @[rob.scala 147:39]
  wire [6:0] _GEN_26421 = io_i_ex_res_packs_1_valid ? _GEN_24245 : _GEN_22069; // @[rob.scala 147:39]
  wire [6:0] _GEN_26422 = io_i_ex_res_packs_1_valid ? _GEN_24246 : _GEN_22070; // @[rob.scala 147:39]
  wire [6:0] _GEN_26423 = io_i_ex_res_packs_1_valid ? _GEN_24247 : _GEN_22071; // @[rob.scala 147:39]
  wire [6:0] _GEN_26424 = io_i_ex_res_packs_1_valid ? _GEN_24248 : _GEN_22072; // @[rob.scala 147:39]
  wire [6:0] _GEN_26425 = io_i_ex_res_packs_1_valid ? _GEN_24249 : _GEN_22073; // @[rob.scala 147:39]
  wire [6:0] _GEN_26426 = io_i_ex_res_packs_1_valid ? _GEN_24250 : _GEN_22074; // @[rob.scala 147:39]
  wire [6:0] _GEN_26427 = io_i_ex_res_packs_1_valid ? _GEN_24251 : _GEN_22075; // @[rob.scala 147:39]
  wire [6:0] _GEN_26428 = io_i_ex_res_packs_1_valid ? _GEN_24252 : _GEN_22076; // @[rob.scala 147:39]
  wire [6:0] _GEN_26429 = io_i_ex_res_packs_1_valid ? _GEN_24253 : _GEN_22077; // @[rob.scala 147:39]
  wire [6:0] _GEN_26430 = io_i_ex_res_packs_1_valid ? _GEN_24254 : _GEN_22078; // @[rob.scala 147:39]
  wire [6:0] _GEN_26431 = io_i_ex_res_packs_1_valid ? _GEN_24255 : _GEN_22079; // @[rob.scala 147:39]
  wire [6:0] _GEN_26432 = io_i_ex_res_packs_1_valid ? _GEN_24256 : _GEN_22080; // @[rob.scala 147:39]
  wire [6:0] _GEN_26433 = io_i_ex_res_packs_1_valid ? _GEN_24257 : _GEN_22081; // @[rob.scala 147:39]
  wire [6:0] _GEN_26434 = io_i_ex_res_packs_1_valid ? _GEN_24258 : _GEN_22082; // @[rob.scala 147:39]
  wire [6:0] _GEN_26435 = io_i_ex_res_packs_1_valid ? _GEN_24259 : _GEN_22083; // @[rob.scala 147:39]
  wire [6:0] _GEN_26436 = io_i_ex_res_packs_1_valid ? _GEN_24260 : _GEN_22084; // @[rob.scala 147:39]
  wire [6:0] _GEN_26437 = io_i_ex_res_packs_1_valid ? _GEN_24261 : _GEN_22085; // @[rob.scala 147:39]
  wire [6:0] _GEN_26438 = io_i_ex_res_packs_1_valid ? _GEN_24262 : _GEN_22086; // @[rob.scala 147:39]
  wire [6:0] _GEN_26439 = io_i_ex_res_packs_1_valid ? _GEN_24263 : _GEN_22087; // @[rob.scala 147:39]
  wire [6:0] _GEN_26440 = io_i_ex_res_packs_1_valid ? _GEN_24264 : _GEN_22088; // @[rob.scala 147:39]
  wire [6:0] _GEN_26441 = io_i_ex_res_packs_1_valid ? _GEN_24265 : _GEN_22089; // @[rob.scala 147:39]
  wire [6:0] _GEN_26442 = io_i_ex_res_packs_1_valid ? _GEN_24266 : _GEN_22090; // @[rob.scala 147:39]
  wire [6:0] _GEN_26443 = io_i_ex_res_packs_1_valid ? _GEN_24267 : _GEN_22091; // @[rob.scala 147:39]
  wire [6:0] _GEN_26444 = io_i_ex_res_packs_1_valid ? _GEN_24268 : _GEN_22092; // @[rob.scala 147:39]
  wire [6:0] _GEN_26445 = io_i_ex_res_packs_1_valid ? _GEN_24269 : _GEN_22093; // @[rob.scala 147:39]
  wire [6:0] _GEN_26446 = io_i_ex_res_packs_1_valid ? _GEN_24270 : _GEN_22094; // @[rob.scala 147:39]
  wire [6:0] _GEN_26447 = io_i_ex_res_packs_1_valid ? _GEN_24271 : _GEN_22095; // @[rob.scala 147:39]
  wire [6:0] _GEN_26448 = io_i_ex_res_packs_1_valid ? _GEN_24272 : _GEN_22096; // @[rob.scala 147:39]
  wire [6:0] _GEN_26449 = io_i_ex_res_packs_1_valid ? _GEN_24273 : _GEN_22097; // @[rob.scala 147:39]
  wire [6:0] _GEN_26450 = io_i_ex_res_packs_1_valid ? _GEN_24274 : _GEN_22098; // @[rob.scala 147:39]
  wire [6:0] _GEN_26451 = io_i_ex_res_packs_1_valid ? _GEN_24275 : _GEN_22099; // @[rob.scala 147:39]
  wire [6:0] _GEN_26452 = io_i_ex_res_packs_1_valid ? _GEN_24276 : _GEN_22100; // @[rob.scala 147:39]
  wire [6:0] _GEN_26453 = io_i_ex_res_packs_1_valid ? _GEN_24277 : _GEN_22101; // @[rob.scala 147:39]
  wire [6:0] _GEN_26454 = io_i_ex_res_packs_1_valid ? _GEN_24278 : _GEN_22102; // @[rob.scala 147:39]
  wire [6:0] _GEN_26455 = io_i_ex_res_packs_1_valid ? _GEN_24279 : _GEN_22103; // @[rob.scala 147:39]
  wire [6:0] _GEN_26456 = io_i_ex_res_packs_1_valid ? _GEN_24280 : _GEN_22104; // @[rob.scala 147:39]
  wire [6:0] _GEN_26457 = io_i_ex_res_packs_1_valid ? _GEN_24281 : _GEN_22105; // @[rob.scala 147:39]
  wire [6:0] _GEN_26458 = io_i_ex_res_packs_1_valid ? _GEN_24282 : _GEN_22106; // @[rob.scala 147:39]
  wire [6:0] _GEN_26459 = io_i_ex_res_packs_1_valid ? _GEN_24283 : _GEN_22107; // @[rob.scala 147:39]
  wire [6:0] _GEN_26460 = io_i_ex_res_packs_1_valid ? _GEN_24284 : _GEN_22108; // @[rob.scala 147:39]
  wire [6:0] _GEN_26461 = io_i_ex_res_packs_1_valid ? _GEN_24285 : _GEN_22109; // @[rob.scala 147:39]
  wire [6:0] _GEN_26462 = io_i_ex_res_packs_1_valid ? _GEN_24286 : _GEN_22110; // @[rob.scala 147:39]
  wire [6:0] _GEN_26463 = io_i_ex_res_packs_1_valid ? _GEN_24287 : _GEN_22111; // @[rob.scala 147:39]
  wire [6:0] _GEN_26464 = io_i_ex_res_packs_1_valid ? _GEN_24288 : _GEN_22112; // @[rob.scala 147:39]
  wire [6:0] _GEN_26465 = io_i_ex_res_packs_1_valid ? _GEN_24289 : _GEN_22113; // @[rob.scala 147:39]
  wire [6:0] _GEN_26466 = io_i_ex_res_packs_1_valid ? _GEN_24290 : _GEN_22114; // @[rob.scala 147:39]
  wire [6:0] _GEN_26467 = io_i_ex_res_packs_1_valid ? _GEN_24291 : _GEN_22115; // @[rob.scala 147:39]
  wire [6:0] _GEN_26468 = io_i_ex_res_packs_1_valid ? _GEN_24292 : _GEN_22116; // @[rob.scala 147:39]
  wire [6:0] _GEN_26469 = io_i_ex_res_packs_1_valid ? _GEN_24293 : _GEN_22117; // @[rob.scala 147:39]
  wire [6:0] _GEN_26470 = io_i_ex_res_packs_1_valid ? _GEN_24294 : _GEN_22118; // @[rob.scala 147:39]
  wire [6:0] _GEN_26471 = io_i_ex_res_packs_1_valid ? _GEN_24295 : _GEN_22119; // @[rob.scala 147:39]
  wire [6:0] _GEN_26472 = io_i_ex_res_packs_1_valid ? _GEN_24296 : _GEN_22120; // @[rob.scala 147:39]
  wire [6:0] _GEN_26473 = io_i_ex_res_packs_1_valid ? _GEN_24297 : _GEN_22121; // @[rob.scala 147:39]
  wire [6:0] _GEN_26474 = io_i_ex_res_packs_1_valid ? _GEN_24298 : _GEN_22122; // @[rob.scala 147:39]
  wire [6:0] _GEN_26475 = io_i_ex_res_packs_1_valid ? _GEN_24299 : _GEN_22123; // @[rob.scala 147:39]
  wire [6:0] _GEN_26476 = io_i_ex_res_packs_1_valid ? _GEN_24300 : _GEN_22124; // @[rob.scala 147:39]
  wire [6:0] _GEN_26477 = io_i_ex_res_packs_1_valid ? _GEN_24301 : _GEN_22125; // @[rob.scala 147:39]
  wire [6:0] _GEN_26478 = io_i_ex_res_packs_1_valid ? _GEN_24302 : _GEN_22126; // @[rob.scala 147:39]
  wire [6:0] _GEN_26479 = io_i_ex_res_packs_1_valid ? _GEN_24303 : _GEN_22127; // @[rob.scala 147:39]
  wire [6:0] _GEN_26480 = io_i_ex_res_packs_1_valid ? _GEN_24304 : _GEN_22128; // @[rob.scala 147:39]
  wire [6:0] _GEN_26481 = io_i_ex_res_packs_1_valid ? _GEN_24305 : _GEN_22129; // @[rob.scala 147:39]
  wire [6:0] _GEN_26482 = io_i_ex_res_packs_1_valid ? _GEN_24306 : _GEN_22130; // @[rob.scala 147:39]
  wire [6:0] _GEN_26483 = io_i_ex_res_packs_1_valid ? _GEN_24307 : _GEN_22131; // @[rob.scala 147:39]
  wire [6:0] _GEN_26484 = io_i_ex_res_packs_1_valid ? _GEN_24308 : _GEN_22132; // @[rob.scala 147:39]
  wire [6:0] _GEN_26485 = io_i_ex_res_packs_1_valid ? _GEN_24309 : _GEN_22133; // @[rob.scala 147:39]
  wire [6:0] _GEN_26486 = io_i_ex_res_packs_1_valid ? _GEN_24310 : _GEN_22134; // @[rob.scala 147:39]
  wire [6:0] _GEN_26487 = io_i_ex_res_packs_1_valid ? _GEN_24311 : _GEN_22135; // @[rob.scala 147:39]
  wire [6:0] _GEN_26488 = io_i_ex_res_packs_1_valid ? _GEN_24312 : _GEN_22136; // @[rob.scala 147:39]
  wire [6:0] _GEN_26489 = io_i_ex_res_packs_1_valid ? _GEN_24313 : _GEN_22137; // @[rob.scala 147:39]
  wire [6:0] _GEN_26490 = io_i_ex_res_packs_1_valid ? _GEN_24314 : _GEN_22138; // @[rob.scala 147:39]
  wire [6:0] _GEN_26491 = io_i_ex_res_packs_1_valid ? _GEN_24315 : _GEN_22139; // @[rob.scala 147:39]
  wire [6:0] _GEN_26492 = io_i_ex_res_packs_1_valid ? _GEN_24316 : _GEN_22140; // @[rob.scala 147:39]
  wire [6:0] _GEN_26493 = io_i_ex_res_packs_1_valid ? _GEN_24317 : _GEN_22141; // @[rob.scala 147:39]
  wire [6:0] _GEN_26494 = io_i_ex_res_packs_1_valid ? _GEN_24318 : _GEN_22142; // @[rob.scala 147:39]
  wire [6:0] _GEN_26495 = io_i_ex_res_packs_1_valid ? _GEN_24319 : _GEN_22143; // @[rob.scala 147:39]
  wire [6:0] _GEN_26496 = io_i_ex_res_packs_1_valid ? _GEN_24320 : _GEN_22144; // @[rob.scala 147:39]
  wire [6:0] _GEN_26497 = io_i_ex_res_packs_1_valid ? _GEN_24321 : _GEN_22145; // @[rob.scala 147:39]
  wire [4:0] _GEN_26498 = io_i_ex_res_packs_1_valid ? _GEN_24322 : _GEN_22146; // @[rob.scala 147:39]
  wire [4:0] _GEN_26499 = io_i_ex_res_packs_1_valid ? _GEN_24323 : _GEN_22147; // @[rob.scala 147:39]
  wire [4:0] _GEN_26500 = io_i_ex_res_packs_1_valid ? _GEN_24324 : _GEN_22148; // @[rob.scala 147:39]
  wire [4:0] _GEN_26501 = io_i_ex_res_packs_1_valid ? _GEN_24325 : _GEN_22149; // @[rob.scala 147:39]
  wire [4:0] _GEN_26502 = io_i_ex_res_packs_1_valid ? _GEN_24326 : _GEN_22150; // @[rob.scala 147:39]
  wire [4:0] _GEN_26503 = io_i_ex_res_packs_1_valid ? _GEN_24327 : _GEN_22151; // @[rob.scala 147:39]
  wire [4:0] _GEN_26504 = io_i_ex_res_packs_1_valid ? _GEN_24328 : _GEN_22152; // @[rob.scala 147:39]
  wire [4:0] _GEN_26505 = io_i_ex_res_packs_1_valid ? _GEN_24329 : _GEN_22153; // @[rob.scala 147:39]
  wire [4:0] _GEN_26506 = io_i_ex_res_packs_1_valid ? _GEN_24330 : _GEN_22154; // @[rob.scala 147:39]
  wire [4:0] _GEN_26507 = io_i_ex_res_packs_1_valid ? _GEN_24331 : _GEN_22155; // @[rob.scala 147:39]
  wire [4:0] _GEN_26508 = io_i_ex_res_packs_1_valid ? _GEN_24332 : _GEN_22156; // @[rob.scala 147:39]
  wire [4:0] _GEN_26509 = io_i_ex_res_packs_1_valid ? _GEN_24333 : _GEN_22157; // @[rob.scala 147:39]
  wire [4:0] _GEN_26510 = io_i_ex_res_packs_1_valid ? _GEN_24334 : _GEN_22158; // @[rob.scala 147:39]
  wire [4:0] _GEN_26511 = io_i_ex_res_packs_1_valid ? _GEN_24335 : _GEN_22159; // @[rob.scala 147:39]
  wire [4:0] _GEN_26512 = io_i_ex_res_packs_1_valid ? _GEN_24336 : _GEN_22160; // @[rob.scala 147:39]
  wire [4:0] _GEN_26513 = io_i_ex_res_packs_1_valid ? _GEN_24337 : _GEN_22161; // @[rob.scala 147:39]
  wire [4:0] _GEN_26514 = io_i_ex_res_packs_1_valid ? _GEN_24338 : _GEN_22162; // @[rob.scala 147:39]
  wire [4:0] _GEN_26515 = io_i_ex_res_packs_1_valid ? _GEN_24339 : _GEN_22163; // @[rob.scala 147:39]
  wire [4:0] _GEN_26516 = io_i_ex_res_packs_1_valid ? _GEN_24340 : _GEN_22164; // @[rob.scala 147:39]
  wire [4:0] _GEN_26517 = io_i_ex_res_packs_1_valid ? _GEN_24341 : _GEN_22165; // @[rob.scala 147:39]
  wire [4:0] _GEN_26518 = io_i_ex_res_packs_1_valid ? _GEN_24342 : _GEN_22166; // @[rob.scala 147:39]
  wire [4:0] _GEN_26519 = io_i_ex_res_packs_1_valid ? _GEN_24343 : _GEN_22167; // @[rob.scala 147:39]
  wire [4:0] _GEN_26520 = io_i_ex_res_packs_1_valid ? _GEN_24344 : _GEN_22168; // @[rob.scala 147:39]
  wire [4:0] _GEN_26521 = io_i_ex_res_packs_1_valid ? _GEN_24345 : _GEN_22169; // @[rob.scala 147:39]
  wire [4:0] _GEN_26522 = io_i_ex_res_packs_1_valid ? _GEN_24346 : _GEN_22170; // @[rob.scala 147:39]
  wire [4:0] _GEN_26523 = io_i_ex_res_packs_1_valid ? _GEN_24347 : _GEN_22171; // @[rob.scala 147:39]
  wire [4:0] _GEN_26524 = io_i_ex_res_packs_1_valid ? _GEN_24348 : _GEN_22172; // @[rob.scala 147:39]
  wire [4:0] _GEN_26525 = io_i_ex_res_packs_1_valid ? _GEN_24349 : _GEN_22173; // @[rob.scala 147:39]
  wire [4:0] _GEN_26526 = io_i_ex_res_packs_1_valid ? _GEN_24350 : _GEN_22174; // @[rob.scala 147:39]
  wire [4:0] _GEN_26527 = io_i_ex_res_packs_1_valid ? _GEN_24351 : _GEN_22175; // @[rob.scala 147:39]
  wire [4:0] _GEN_26528 = io_i_ex_res_packs_1_valid ? _GEN_24352 : _GEN_22176; // @[rob.scala 147:39]
  wire [4:0] _GEN_26529 = io_i_ex_res_packs_1_valid ? _GEN_24353 : _GEN_22177; // @[rob.scala 147:39]
  wire [4:0] _GEN_26530 = io_i_ex_res_packs_1_valid ? _GEN_24354 : _GEN_22178; // @[rob.scala 147:39]
  wire [4:0] _GEN_26531 = io_i_ex_res_packs_1_valid ? _GEN_24355 : _GEN_22179; // @[rob.scala 147:39]
  wire [4:0] _GEN_26532 = io_i_ex_res_packs_1_valid ? _GEN_24356 : _GEN_22180; // @[rob.scala 147:39]
  wire [4:0] _GEN_26533 = io_i_ex_res_packs_1_valid ? _GEN_24357 : _GEN_22181; // @[rob.scala 147:39]
  wire [4:0] _GEN_26534 = io_i_ex_res_packs_1_valid ? _GEN_24358 : _GEN_22182; // @[rob.scala 147:39]
  wire [4:0] _GEN_26535 = io_i_ex_res_packs_1_valid ? _GEN_24359 : _GEN_22183; // @[rob.scala 147:39]
  wire [4:0] _GEN_26536 = io_i_ex_res_packs_1_valid ? _GEN_24360 : _GEN_22184; // @[rob.scala 147:39]
  wire [4:0] _GEN_26537 = io_i_ex_res_packs_1_valid ? _GEN_24361 : _GEN_22185; // @[rob.scala 147:39]
  wire [4:0] _GEN_26538 = io_i_ex_res_packs_1_valid ? _GEN_24362 : _GEN_22186; // @[rob.scala 147:39]
  wire [4:0] _GEN_26539 = io_i_ex_res_packs_1_valid ? _GEN_24363 : _GEN_22187; // @[rob.scala 147:39]
  wire [4:0] _GEN_26540 = io_i_ex_res_packs_1_valid ? _GEN_24364 : _GEN_22188; // @[rob.scala 147:39]
  wire [4:0] _GEN_26541 = io_i_ex_res_packs_1_valid ? _GEN_24365 : _GEN_22189; // @[rob.scala 147:39]
  wire [4:0] _GEN_26542 = io_i_ex_res_packs_1_valid ? _GEN_24366 : _GEN_22190; // @[rob.scala 147:39]
  wire [4:0] _GEN_26543 = io_i_ex_res_packs_1_valid ? _GEN_24367 : _GEN_22191; // @[rob.scala 147:39]
  wire [4:0] _GEN_26544 = io_i_ex_res_packs_1_valid ? _GEN_24368 : _GEN_22192; // @[rob.scala 147:39]
  wire [4:0] _GEN_26545 = io_i_ex_res_packs_1_valid ? _GEN_24369 : _GEN_22193; // @[rob.scala 147:39]
  wire [4:0] _GEN_26546 = io_i_ex_res_packs_1_valid ? _GEN_24370 : _GEN_22194; // @[rob.scala 147:39]
  wire [4:0] _GEN_26547 = io_i_ex_res_packs_1_valid ? _GEN_24371 : _GEN_22195; // @[rob.scala 147:39]
  wire [4:0] _GEN_26548 = io_i_ex_res_packs_1_valid ? _GEN_24372 : _GEN_22196; // @[rob.scala 147:39]
  wire [4:0] _GEN_26549 = io_i_ex_res_packs_1_valid ? _GEN_24373 : _GEN_22197; // @[rob.scala 147:39]
  wire [4:0] _GEN_26550 = io_i_ex_res_packs_1_valid ? _GEN_24374 : _GEN_22198; // @[rob.scala 147:39]
  wire [4:0] _GEN_26551 = io_i_ex_res_packs_1_valid ? _GEN_24375 : _GEN_22199; // @[rob.scala 147:39]
  wire [4:0] _GEN_26552 = io_i_ex_res_packs_1_valid ? _GEN_24376 : _GEN_22200; // @[rob.scala 147:39]
  wire [4:0] _GEN_26553 = io_i_ex_res_packs_1_valid ? _GEN_24377 : _GEN_22201; // @[rob.scala 147:39]
  wire [4:0] _GEN_26554 = io_i_ex_res_packs_1_valid ? _GEN_24378 : _GEN_22202; // @[rob.scala 147:39]
  wire [4:0] _GEN_26555 = io_i_ex_res_packs_1_valid ? _GEN_24379 : _GEN_22203; // @[rob.scala 147:39]
  wire [4:0] _GEN_26556 = io_i_ex_res_packs_1_valid ? _GEN_24380 : _GEN_22204; // @[rob.scala 147:39]
  wire [4:0] _GEN_26557 = io_i_ex_res_packs_1_valid ? _GEN_24381 : _GEN_22205; // @[rob.scala 147:39]
  wire [4:0] _GEN_26558 = io_i_ex_res_packs_1_valid ? _GEN_24382 : _GEN_22206; // @[rob.scala 147:39]
  wire [4:0] _GEN_26559 = io_i_ex_res_packs_1_valid ? _GEN_24383 : _GEN_22207; // @[rob.scala 147:39]
  wire [4:0] _GEN_26560 = io_i_ex_res_packs_1_valid ? _GEN_24384 : _GEN_22208; // @[rob.scala 147:39]
  wire [4:0] _GEN_26561 = io_i_ex_res_packs_1_valid ? _GEN_24385 : _GEN_22209; // @[rob.scala 147:39]
  wire [63:0] _GEN_27202 = io_i_ex_res_packs_1_valid ? _GEN_25026 : _GEN_22850; // @[rob.scala 147:39]
  wire [63:0] _GEN_27203 = io_i_ex_res_packs_1_valid ? _GEN_25027 : _GEN_22851; // @[rob.scala 147:39]
  wire [63:0] _GEN_27204 = io_i_ex_res_packs_1_valid ? _GEN_25028 : _GEN_22852; // @[rob.scala 147:39]
  wire [63:0] _GEN_27205 = io_i_ex_res_packs_1_valid ? _GEN_25029 : _GEN_22853; // @[rob.scala 147:39]
  wire [63:0] _GEN_27206 = io_i_ex_res_packs_1_valid ? _GEN_25030 : _GEN_22854; // @[rob.scala 147:39]
  wire [63:0] _GEN_27207 = io_i_ex_res_packs_1_valid ? _GEN_25031 : _GEN_22855; // @[rob.scala 147:39]
  wire [63:0] _GEN_27208 = io_i_ex_res_packs_1_valid ? _GEN_25032 : _GEN_22856; // @[rob.scala 147:39]
  wire [63:0] _GEN_27209 = io_i_ex_res_packs_1_valid ? _GEN_25033 : _GEN_22857; // @[rob.scala 147:39]
  wire [63:0] _GEN_27210 = io_i_ex_res_packs_1_valid ? _GEN_25034 : _GEN_22858; // @[rob.scala 147:39]
  wire [63:0] _GEN_27211 = io_i_ex_res_packs_1_valid ? _GEN_25035 : _GEN_22859; // @[rob.scala 147:39]
  wire [63:0] _GEN_27212 = io_i_ex_res_packs_1_valid ? _GEN_25036 : _GEN_22860; // @[rob.scala 147:39]
  wire [63:0] _GEN_27213 = io_i_ex_res_packs_1_valid ? _GEN_25037 : _GEN_22861; // @[rob.scala 147:39]
  wire [63:0] _GEN_27214 = io_i_ex_res_packs_1_valid ? _GEN_25038 : _GEN_22862; // @[rob.scala 147:39]
  wire [63:0] _GEN_27215 = io_i_ex_res_packs_1_valid ? _GEN_25039 : _GEN_22863; // @[rob.scala 147:39]
  wire [63:0] _GEN_27216 = io_i_ex_res_packs_1_valid ? _GEN_25040 : _GEN_22864; // @[rob.scala 147:39]
  wire [63:0] _GEN_27217 = io_i_ex_res_packs_1_valid ? _GEN_25041 : _GEN_22865; // @[rob.scala 147:39]
  wire [63:0] _GEN_27218 = io_i_ex_res_packs_1_valid ? _GEN_25042 : _GEN_22866; // @[rob.scala 147:39]
  wire [63:0] _GEN_27219 = io_i_ex_res_packs_1_valid ? _GEN_25043 : _GEN_22867; // @[rob.scala 147:39]
  wire [63:0] _GEN_27220 = io_i_ex_res_packs_1_valid ? _GEN_25044 : _GEN_22868; // @[rob.scala 147:39]
  wire [63:0] _GEN_27221 = io_i_ex_res_packs_1_valid ? _GEN_25045 : _GEN_22869; // @[rob.scala 147:39]
  wire [63:0] _GEN_27222 = io_i_ex_res_packs_1_valid ? _GEN_25046 : _GEN_22870; // @[rob.scala 147:39]
  wire [63:0] _GEN_27223 = io_i_ex_res_packs_1_valid ? _GEN_25047 : _GEN_22871; // @[rob.scala 147:39]
  wire [63:0] _GEN_27224 = io_i_ex_res_packs_1_valid ? _GEN_25048 : _GEN_22872; // @[rob.scala 147:39]
  wire [63:0] _GEN_27225 = io_i_ex_res_packs_1_valid ? _GEN_25049 : _GEN_22873; // @[rob.scala 147:39]
  wire [63:0] _GEN_27226 = io_i_ex_res_packs_1_valid ? _GEN_25050 : _GEN_22874; // @[rob.scala 147:39]
  wire [63:0] _GEN_27227 = io_i_ex_res_packs_1_valid ? _GEN_25051 : _GEN_22875; // @[rob.scala 147:39]
  wire [63:0] _GEN_27228 = io_i_ex_res_packs_1_valid ? _GEN_25052 : _GEN_22876; // @[rob.scala 147:39]
  wire [63:0] _GEN_27229 = io_i_ex_res_packs_1_valid ? _GEN_25053 : _GEN_22877; // @[rob.scala 147:39]
  wire [63:0] _GEN_27230 = io_i_ex_res_packs_1_valid ? _GEN_25054 : _GEN_22878; // @[rob.scala 147:39]
  wire [63:0] _GEN_27231 = io_i_ex_res_packs_1_valid ? _GEN_25055 : _GEN_22879; // @[rob.scala 147:39]
  wire [63:0] _GEN_27232 = io_i_ex_res_packs_1_valid ? _GEN_25056 : _GEN_22880; // @[rob.scala 147:39]
  wire [63:0] _GEN_27233 = io_i_ex_res_packs_1_valid ? _GEN_25057 : _GEN_22881; // @[rob.scala 147:39]
  wire [63:0] _GEN_27234 = io_i_ex_res_packs_1_valid ? _GEN_25058 : _GEN_22882; // @[rob.scala 147:39]
  wire [63:0] _GEN_27235 = io_i_ex_res_packs_1_valid ? _GEN_25059 : _GEN_22883; // @[rob.scala 147:39]
  wire [63:0] _GEN_27236 = io_i_ex_res_packs_1_valid ? _GEN_25060 : _GEN_22884; // @[rob.scala 147:39]
  wire [63:0] _GEN_27237 = io_i_ex_res_packs_1_valid ? _GEN_25061 : _GEN_22885; // @[rob.scala 147:39]
  wire [63:0] _GEN_27238 = io_i_ex_res_packs_1_valid ? _GEN_25062 : _GEN_22886; // @[rob.scala 147:39]
  wire [63:0] _GEN_27239 = io_i_ex_res_packs_1_valid ? _GEN_25063 : _GEN_22887; // @[rob.scala 147:39]
  wire [63:0] _GEN_27240 = io_i_ex_res_packs_1_valid ? _GEN_25064 : _GEN_22888; // @[rob.scala 147:39]
  wire [63:0] _GEN_27241 = io_i_ex_res_packs_1_valid ? _GEN_25065 : _GEN_22889; // @[rob.scala 147:39]
  wire [63:0] _GEN_27242 = io_i_ex_res_packs_1_valid ? _GEN_25066 : _GEN_22890; // @[rob.scala 147:39]
  wire [63:0] _GEN_27243 = io_i_ex_res_packs_1_valid ? _GEN_25067 : _GEN_22891; // @[rob.scala 147:39]
  wire [63:0] _GEN_27244 = io_i_ex_res_packs_1_valid ? _GEN_25068 : _GEN_22892; // @[rob.scala 147:39]
  wire [63:0] _GEN_27245 = io_i_ex_res_packs_1_valid ? _GEN_25069 : _GEN_22893; // @[rob.scala 147:39]
  wire [63:0] _GEN_27246 = io_i_ex_res_packs_1_valid ? _GEN_25070 : _GEN_22894; // @[rob.scala 147:39]
  wire [63:0] _GEN_27247 = io_i_ex_res_packs_1_valid ? _GEN_25071 : _GEN_22895; // @[rob.scala 147:39]
  wire [63:0] _GEN_27248 = io_i_ex_res_packs_1_valid ? _GEN_25072 : _GEN_22896; // @[rob.scala 147:39]
  wire [63:0] _GEN_27249 = io_i_ex_res_packs_1_valid ? _GEN_25073 : _GEN_22897; // @[rob.scala 147:39]
  wire [63:0] _GEN_27250 = io_i_ex_res_packs_1_valid ? _GEN_25074 : _GEN_22898; // @[rob.scala 147:39]
  wire [63:0] _GEN_27251 = io_i_ex_res_packs_1_valid ? _GEN_25075 : _GEN_22899; // @[rob.scala 147:39]
  wire [63:0] _GEN_27252 = io_i_ex_res_packs_1_valid ? _GEN_25076 : _GEN_22900; // @[rob.scala 147:39]
  wire [63:0] _GEN_27253 = io_i_ex_res_packs_1_valid ? _GEN_25077 : _GEN_22901; // @[rob.scala 147:39]
  wire [63:0] _GEN_27254 = io_i_ex_res_packs_1_valid ? _GEN_25078 : _GEN_22902; // @[rob.scala 147:39]
  wire [63:0] _GEN_27255 = io_i_ex_res_packs_1_valid ? _GEN_25079 : _GEN_22903; // @[rob.scala 147:39]
  wire [63:0] _GEN_27256 = io_i_ex_res_packs_1_valid ? _GEN_25080 : _GEN_22904; // @[rob.scala 147:39]
  wire [63:0] _GEN_27257 = io_i_ex_res_packs_1_valid ? _GEN_25081 : _GEN_22905; // @[rob.scala 147:39]
  wire [63:0] _GEN_27258 = io_i_ex_res_packs_1_valid ? _GEN_25082 : _GEN_22906; // @[rob.scala 147:39]
  wire [63:0] _GEN_27259 = io_i_ex_res_packs_1_valid ? _GEN_25083 : _GEN_22907; // @[rob.scala 147:39]
  wire [63:0] _GEN_27260 = io_i_ex_res_packs_1_valid ? _GEN_25084 : _GEN_22908; // @[rob.scala 147:39]
  wire [63:0] _GEN_27261 = io_i_ex_res_packs_1_valid ? _GEN_25085 : _GEN_22909; // @[rob.scala 147:39]
  wire [63:0] _GEN_27262 = io_i_ex_res_packs_1_valid ? _GEN_25086 : _GEN_22910; // @[rob.scala 147:39]
  wire [63:0] _GEN_27263 = io_i_ex_res_packs_1_valid ? _GEN_25087 : _GEN_22911; // @[rob.scala 147:39]
  wire [63:0] _GEN_27264 = io_i_ex_res_packs_1_valid ? _GEN_25088 : _GEN_22912; // @[rob.scala 147:39]
  wire [63:0] _GEN_27265 = io_i_ex_res_packs_1_valid ? _GEN_25089 : _GEN_22913; // @[rob.scala 147:39]
  wire [63:0] _GEN_27266 = io_i_ex_res_packs_1_valid ? _GEN_25090 : _GEN_22914; // @[rob.scala 147:39]
  wire [63:0] _GEN_27267 = io_i_ex_res_packs_1_valid ? _GEN_25091 : _GEN_22915; // @[rob.scala 147:39]
  wire [63:0] _GEN_27268 = io_i_ex_res_packs_1_valid ? _GEN_25092 : _GEN_22916; // @[rob.scala 147:39]
  wire [63:0] _GEN_27269 = io_i_ex_res_packs_1_valid ? _GEN_25093 : _GEN_22917; // @[rob.scala 147:39]
  wire [63:0] _GEN_27270 = io_i_ex_res_packs_1_valid ? _GEN_25094 : _GEN_22918; // @[rob.scala 147:39]
  wire [63:0] _GEN_27271 = io_i_ex_res_packs_1_valid ? _GEN_25095 : _GEN_22919; // @[rob.scala 147:39]
  wire [63:0] _GEN_27272 = io_i_ex_res_packs_1_valid ? _GEN_25096 : _GEN_22920; // @[rob.scala 147:39]
  wire [63:0] _GEN_27273 = io_i_ex_res_packs_1_valid ? _GEN_25097 : _GEN_22921; // @[rob.scala 147:39]
  wire [63:0] _GEN_27274 = io_i_ex_res_packs_1_valid ? _GEN_25098 : _GEN_22922; // @[rob.scala 147:39]
  wire [63:0] _GEN_27275 = io_i_ex_res_packs_1_valid ? _GEN_25099 : _GEN_22923; // @[rob.scala 147:39]
  wire [63:0] _GEN_27276 = io_i_ex_res_packs_1_valid ? _GEN_25100 : _GEN_22924; // @[rob.scala 147:39]
  wire [63:0] _GEN_27277 = io_i_ex_res_packs_1_valid ? _GEN_25101 : _GEN_22925; // @[rob.scala 147:39]
  wire [63:0] _GEN_27278 = io_i_ex_res_packs_1_valid ? _GEN_25102 : _GEN_22926; // @[rob.scala 147:39]
  wire [63:0] _GEN_27279 = io_i_ex_res_packs_1_valid ? _GEN_25103 : _GEN_22927; // @[rob.scala 147:39]
  wire [63:0] _GEN_27280 = io_i_ex_res_packs_1_valid ? _GEN_25104 : _GEN_22928; // @[rob.scala 147:39]
  wire [63:0] _GEN_27281 = io_i_ex_res_packs_1_valid ? _GEN_25105 : _GEN_22929; // @[rob.scala 147:39]
  wire [63:0] _GEN_27282 = io_i_ex_res_packs_1_valid ? _GEN_25106 : _GEN_22930; // @[rob.scala 147:39]
  wire [63:0] _GEN_27283 = io_i_ex_res_packs_1_valid ? _GEN_25107 : _GEN_22931; // @[rob.scala 147:39]
  wire [63:0] _GEN_27284 = io_i_ex_res_packs_1_valid ? _GEN_25108 : _GEN_22932; // @[rob.scala 147:39]
  wire [63:0] _GEN_27285 = io_i_ex_res_packs_1_valid ? _GEN_25109 : _GEN_22933; // @[rob.scala 147:39]
  wire [63:0] _GEN_27286 = io_i_ex_res_packs_1_valid ? _GEN_25110 : _GEN_22934; // @[rob.scala 147:39]
  wire [63:0] _GEN_27287 = io_i_ex_res_packs_1_valid ? _GEN_25111 : _GEN_22935; // @[rob.scala 147:39]
  wire [63:0] _GEN_27288 = io_i_ex_res_packs_1_valid ? _GEN_25112 : _GEN_22936; // @[rob.scala 147:39]
  wire [63:0] _GEN_27289 = io_i_ex_res_packs_1_valid ? _GEN_25113 : _GEN_22937; // @[rob.scala 147:39]
  wire [63:0] _GEN_27290 = io_i_ex_res_packs_1_valid ? _GEN_25114 : _GEN_22938; // @[rob.scala 147:39]
  wire [63:0] _GEN_27291 = io_i_ex_res_packs_1_valid ? _GEN_25115 : _GEN_22939; // @[rob.scala 147:39]
  wire [63:0] _GEN_27292 = io_i_ex_res_packs_1_valid ? _GEN_25116 : _GEN_22940; // @[rob.scala 147:39]
  wire [63:0] _GEN_27293 = io_i_ex_res_packs_1_valid ? _GEN_25117 : _GEN_22941; // @[rob.scala 147:39]
  wire [63:0] _GEN_27294 = io_i_ex_res_packs_1_valid ? _GEN_25118 : _GEN_22942; // @[rob.scala 147:39]
  wire [63:0] _GEN_27295 = io_i_ex_res_packs_1_valid ? _GEN_25119 : _GEN_22943; // @[rob.scala 147:39]
  wire [63:0] _GEN_27296 = io_i_ex_res_packs_1_valid ? _GEN_25120 : _GEN_22944; // @[rob.scala 147:39]
  wire [63:0] _GEN_27297 = io_i_ex_res_packs_1_valid ? _GEN_25121 : _GEN_22945; // @[rob.scala 147:39]
  wire [63:0] _GEN_27298 = io_i_ex_res_packs_1_valid ? _GEN_25122 : _GEN_22946; // @[rob.scala 147:39]
  wire [63:0] _GEN_27299 = io_i_ex_res_packs_1_valid ? _GEN_25123 : _GEN_22947; // @[rob.scala 147:39]
  wire [63:0] _GEN_27300 = io_i_ex_res_packs_1_valid ? _GEN_25124 : _GEN_22948; // @[rob.scala 147:39]
  wire [63:0] _GEN_27301 = io_i_ex_res_packs_1_valid ? _GEN_25125 : _GEN_22949; // @[rob.scala 147:39]
  wire [63:0] _GEN_27302 = io_i_ex_res_packs_1_valid ? _GEN_25126 : _GEN_22950; // @[rob.scala 147:39]
  wire [63:0] _GEN_27303 = io_i_ex_res_packs_1_valid ? _GEN_25127 : _GEN_22951; // @[rob.scala 147:39]
  wire [63:0] _GEN_27304 = io_i_ex_res_packs_1_valid ? _GEN_25128 : _GEN_22952; // @[rob.scala 147:39]
  wire [63:0] _GEN_27305 = io_i_ex_res_packs_1_valid ? _GEN_25129 : _GEN_22953; // @[rob.scala 147:39]
  wire [63:0] _GEN_27306 = io_i_ex_res_packs_1_valid ? _GEN_25130 : _GEN_22954; // @[rob.scala 147:39]
  wire [63:0] _GEN_27307 = io_i_ex_res_packs_1_valid ? _GEN_25131 : _GEN_22955; // @[rob.scala 147:39]
  wire [63:0] _GEN_27308 = io_i_ex_res_packs_1_valid ? _GEN_25132 : _GEN_22956; // @[rob.scala 147:39]
  wire [63:0] _GEN_27309 = io_i_ex_res_packs_1_valid ? _GEN_25133 : _GEN_22957; // @[rob.scala 147:39]
  wire [63:0] _GEN_27310 = io_i_ex_res_packs_1_valid ? _GEN_25134 : _GEN_22958; // @[rob.scala 147:39]
  wire [63:0] _GEN_27311 = io_i_ex_res_packs_1_valid ? _GEN_25135 : _GEN_22959; // @[rob.scala 147:39]
  wire [63:0] _GEN_27312 = io_i_ex_res_packs_1_valid ? _GEN_25136 : _GEN_22960; // @[rob.scala 147:39]
  wire [63:0] _GEN_27313 = io_i_ex_res_packs_1_valid ? _GEN_25137 : _GEN_22961; // @[rob.scala 147:39]
  wire [63:0] _GEN_27314 = io_i_ex_res_packs_1_valid ? _GEN_25138 : _GEN_22962; // @[rob.scala 147:39]
  wire [63:0] _GEN_27315 = io_i_ex_res_packs_1_valid ? _GEN_25139 : _GEN_22963; // @[rob.scala 147:39]
  wire [63:0] _GEN_27316 = io_i_ex_res_packs_1_valid ? _GEN_25140 : _GEN_22964; // @[rob.scala 147:39]
  wire [63:0] _GEN_27317 = io_i_ex_res_packs_1_valid ? _GEN_25141 : _GEN_22965; // @[rob.scala 147:39]
  wire [63:0] _GEN_27318 = io_i_ex_res_packs_1_valid ? _GEN_25142 : _GEN_22966; // @[rob.scala 147:39]
  wire [63:0] _GEN_27319 = io_i_ex_res_packs_1_valid ? _GEN_25143 : _GEN_22967; // @[rob.scala 147:39]
  wire [63:0] _GEN_27320 = io_i_ex_res_packs_1_valid ? _GEN_25144 : _GEN_22968; // @[rob.scala 147:39]
  wire [63:0] _GEN_27321 = io_i_ex_res_packs_1_valid ? _GEN_25145 : _GEN_22969; // @[rob.scala 147:39]
  wire [63:0] _GEN_27322 = io_i_ex_res_packs_1_valid ? _GEN_25146 : _GEN_22970; // @[rob.scala 147:39]
  wire [63:0] _GEN_27323 = io_i_ex_res_packs_1_valid ? _GEN_25147 : _GEN_22971; // @[rob.scala 147:39]
  wire [63:0] _GEN_27324 = io_i_ex_res_packs_1_valid ? _GEN_25148 : _GEN_22972; // @[rob.scala 147:39]
  wire [63:0] _GEN_27325 = io_i_ex_res_packs_1_valid ? _GEN_25149 : _GEN_22973; // @[rob.scala 147:39]
  wire [63:0] _GEN_27326 = io_i_ex_res_packs_1_valid ? _GEN_25150 : _GEN_22974; // @[rob.scala 147:39]
  wire [63:0] _GEN_27327 = io_i_ex_res_packs_1_valid ? _GEN_25151 : _GEN_22975; // @[rob.scala 147:39]
  wire [63:0] _GEN_27328 = io_i_ex_res_packs_1_valid ? _GEN_25152 : _GEN_22976; // @[rob.scala 147:39]
  wire [63:0] _GEN_27329 = io_i_ex_res_packs_1_valid ? _GEN_25153 : _GEN_22977; // @[rob.scala 147:39]
  wire [4:0] _GEN_27586 = io_i_ex_res_packs_1_valid ? _GEN_25410 : _GEN_23234; // @[rob.scala 147:39]
  wire [4:0] _GEN_27587 = io_i_ex_res_packs_1_valid ? _GEN_25411 : _GEN_23235; // @[rob.scala 147:39]
  wire [4:0] _GEN_27588 = io_i_ex_res_packs_1_valid ? _GEN_25412 : _GEN_23236; // @[rob.scala 147:39]
  wire [4:0] _GEN_27589 = io_i_ex_res_packs_1_valid ? _GEN_25413 : _GEN_23237; // @[rob.scala 147:39]
  wire [4:0] _GEN_27590 = io_i_ex_res_packs_1_valid ? _GEN_25414 : _GEN_23238; // @[rob.scala 147:39]
  wire [4:0] _GEN_27591 = io_i_ex_res_packs_1_valid ? _GEN_25415 : _GEN_23239; // @[rob.scala 147:39]
  wire [4:0] _GEN_27592 = io_i_ex_res_packs_1_valid ? _GEN_25416 : _GEN_23240; // @[rob.scala 147:39]
  wire [4:0] _GEN_27593 = io_i_ex_res_packs_1_valid ? _GEN_25417 : _GEN_23241; // @[rob.scala 147:39]
  wire [4:0] _GEN_27594 = io_i_ex_res_packs_1_valid ? _GEN_25418 : _GEN_23242; // @[rob.scala 147:39]
  wire [4:0] _GEN_27595 = io_i_ex_res_packs_1_valid ? _GEN_25419 : _GEN_23243; // @[rob.scala 147:39]
  wire [4:0] _GEN_27596 = io_i_ex_res_packs_1_valid ? _GEN_25420 : _GEN_23244; // @[rob.scala 147:39]
  wire [4:0] _GEN_27597 = io_i_ex_res_packs_1_valid ? _GEN_25421 : _GEN_23245; // @[rob.scala 147:39]
  wire [4:0] _GEN_27598 = io_i_ex_res_packs_1_valid ? _GEN_25422 : _GEN_23246; // @[rob.scala 147:39]
  wire [4:0] _GEN_27599 = io_i_ex_res_packs_1_valid ? _GEN_25423 : _GEN_23247; // @[rob.scala 147:39]
  wire [4:0] _GEN_27600 = io_i_ex_res_packs_1_valid ? _GEN_25424 : _GEN_23248; // @[rob.scala 147:39]
  wire [4:0] _GEN_27601 = io_i_ex_res_packs_1_valid ? _GEN_25425 : _GEN_23249; // @[rob.scala 147:39]
  wire [4:0] _GEN_27602 = io_i_ex_res_packs_1_valid ? _GEN_25426 : _GEN_23250; // @[rob.scala 147:39]
  wire [4:0] _GEN_27603 = io_i_ex_res_packs_1_valid ? _GEN_25427 : _GEN_23251; // @[rob.scala 147:39]
  wire [4:0] _GEN_27604 = io_i_ex_res_packs_1_valid ? _GEN_25428 : _GEN_23252; // @[rob.scala 147:39]
  wire [4:0] _GEN_27605 = io_i_ex_res_packs_1_valid ? _GEN_25429 : _GEN_23253; // @[rob.scala 147:39]
  wire [4:0] _GEN_27606 = io_i_ex_res_packs_1_valid ? _GEN_25430 : _GEN_23254; // @[rob.scala 147:39]
  wire [4:0] _GEN_27607 = io_i_ex_res_packs_1_valid ? _GEN_25431 : _GEN_23255; // @[rob.scala 147:39]
  wire [4:0] _GEN_27608 = io_i_ex_res_packs_1_valid ? _GEN_25432 : _GEN_23256; // @[rob.scala 147:39]
  wire [4:0] _GEN_27609 = io_i_ex_res_packs_1_valid ? _GEN_25433 : _GEN_23257; // @[rob.scala 147:39]
  wire [4:0] _GEN_27610 = io_i_ex_res_packs_1_valid ? _GEN_25434 : _GEN_23258; // @[rob.scala 147:39]
  wire [4:0] _GEN_27611 = io_i_ex_res_packs_1_valid ? _GEN_25435 : _GEN_23259; // @[rob.scala 147:39]
  wire [4:0] _GEN_27612 = io_i_ex_res_packs_1_valid ? _GEN_25436 : _GEN_23260; // @[rob.scala 147:39]
  wire [4:0] _GEN_27613 = io_i_ex_res_packs_1_valid ? _GEN_25437 : _GEN_23261; // @[rob.scala 147:39]
  wire [4:0] _GEN_27614 = io_i_ex_res_packs_1_valid ? _GEN_25438 : _GEN_23262; // @[rob.scala 147:39]
  wire [4:0] _GEN_27615 = io_i_ex_res_packs_1_valid ? _GEN_25439 : _GEN_23263; // @[rob.scala 147:39]
  wire [4:0] _GEN_27616 = io_i_ex_res_packs_1_valid ? _GEN_25440 : _GEN_23264; // @[rob.scala 147:39]
  wire [4:0] _GEN_27617 = io_i_ex_res_packs_1_valid ? _GEN_25441 : _GEN_23265; // @[rob.scala 147:39]
  wire [4:0] _GEN_27618 = io_i_ex_res_packs_1_valid ? _GEN_25442 : _GEN_23266; // @[rob.scala 147:39]
  wire [4:0] _GEN_27619 = io_i_ex_res_packs_1_valid ? _GEN_25443 : _GEN_23267; // @[rob.scala 147:39]
  wire [4:0] _GEN_27620 = io_i_ex_res_packs_1_valid ? _GEN_25444 : _GEN_23268; // @[rob.scala 147:39]
  wire [4:0] _GEN_27621 = io_i_ex_res_packs_1_valid ? _GEN_25445 : _GEN_23269; // @[rob.scala 147:39]
  wire [4:0] _GEN_27622 = io_i_ex_res_packs_1_valid ? _GEN_25446 : _GEN_23270; // @[rob.scala 147:39]
  wire [4:0] _GEN_27623 = io_i_ex_res_packs_1_valid ? _GEN_25447 : _GEN_23271; // @[rob.scala 147:39]
  wire [4:0] _GEN_27624 = io_i_ex_res_packs_1_valid ? _GEN_25448 : _GEN_23272; // @[rob.scala 147:39]
  wire [4:0] _GEN_27625 = io_i_ex_res_packs_1_valid ? _GEN_25449 : _GEN_23273; // @[rob.scala 147:39]
  wire [4:0] _GEN_27626 = io_i_ex_res_packs_1_valid ? _GEN_25450 : _GEN_23274; // @[rob.scala 147:39]
  wire [4:0] _GEN_27627 = io_i_ex_res_packs_1_valid ? _GEN_25451 : _GEN_23275; // @[rob.scala 147:39]
  wire [4:0] _GEN_27628 = io_i_ex_res_packs_1_valid ? _GEN_25452 : _GEN_23276; // @[rob.scala 147:39]
  wire [4:0] _GEN_27629 = io_i_ex_res_packs_1_valid ? _GEN_25453 : _GEN_23277; // @[rob.scala 147:39]
  wire [4:0] _GEN_27630 = io_i_ex_res_packs_1_valid ? _GEN_25454 : _GEN_23278; // @[rob.scala 147:39]
  wire [4:0] _GEN_27631 = io_i_ex_res_packs_1_valid ? _GEN_25455 : _GEN_23279; // @[rob.scala 147:39]
  wire [4:0] _GEN_27632 = io_i_ex_res_packs_1_valid ? _GEN_25456 : _GEN_23280; // @[rob.scala 147:39]
  wire [4:0] _GEN_27633 = io_i_ex_res_packs_1_valid ? _GEN_25457 : _GEN_23281; // @[rob.scala 147:39]
  wire [4:0] _GEN_27634 = io_i_ex_res_packs_1_valid ? _GEN_25458 : _GEN_23282; // @[rob.scala 147:39]
  wire [4:0] _GEN_27635 = io_i_ex_res_packs_1_valid ? _GEN_25459 : _GEN_23283; // @[rob.scala 147:39]
  wire [4:0] _GEN_27636 = io_i_ex_res_packs_1_valid ? _GEN_25460 : _GEN_23284; // @[rob.scala 147:39]
  wire [4:0] _GEN_27637 = io_i_ex_res_packs_1_valid ? _GEN_25461 : _GEN_23285; // @[rob.scala 147:39]
  wire [4:0] _GEN_27638 = io_i_ex_res_packs_1_valid ? _GEN_25462 : _GEN_23286; // @[rob.scala 147:39]
  wire [4:0] _GEN_27639 = io_i_ex_res_packs_1_valid ? _GEN_25463 : _GEN_23287; // @[rob.scala 147:39]
  wire [4:0] _GEN_27640 = io_i_ex_res_packs_1_valid ? _GEN_25464 : _GEN_23288; // @[rob.scala 147:39]
  wire [4:0] _GEN_27641 = io_i_ex_res_packs_1_valid ? _GEN_25465 : _GEN_23289; // @[rob.scala 147:39]
  wire [4:0] _GEN_27642 = io_i_ex_res_packs_1_valid ? _GEN_25466 : _GEN_23290; // @[rob.scala 147:39]
  wire [4:0] _GEN_27643 = io_i_ex_res_packs_1_valid ? _GEN_25467 : _GEN_23291; // @[rob.scala 147:39]
  wire [4:0] _GEN_27644 = io_i_ex_res_packs_1_valid ? _GEN_25468 : _GEN_23292; // @[rob.scala 147:39]
  wire [4:0] _GEN_27645 = io_i_ex_res_packs_1_valid ? _GEN_25469 : _GEN_23293; // @[rob.scala 147:39]
  wire [4:0] _GEN_27646 = io_i_ex_res_packs_1_valid ? _GEN_25470 : _GEN_23294; // @[rob.scala 147:39]
  wire [4:0] _GEN_27647 = io_i_ex_res_packs_1_valid ? _GEN_25471 : _GEN_23295; // @[rob.scala 147:39]
  wire [4:0] _GEN_27648 = io_i_ex_res_packs_1_valid ? _GEN_25472 : _GEN_23296; // @[rob.scala 147:39]
  wire [4:0] _GEN_27649 = io_i_ex_res_packs_1_valid ? _GEN_25473 : _GEN_23297; // @[rob.scala 147:39]
  wire  _GEN_27842 = io_i_ex_res_packs_1_valid ? _GEN_25666 : _GEN_23490; // @[rob.scala 147:39]
  wire  _GEN_27843 = io_i_ex_res_packs_1_valid ? _GEN_25667 : _GEN_23491; // @[rob.scala 147:39]
  wire  _GEN_27844 = io_i_ex_res_packs_1_valid ? _GEN_25668 : _GEN_23492; // @[rob.scala 147:39]
  wire  _GEN_27845 = io_i_ex_res_packs_1_valid ? _GEN_25669 : _GEN_23493; // @[rob.scala 147:39]
  wire  _GEN_27846 = io_i_ex_res_packs_1_valid ? _GEN_25670 : _GEN_23494; // @[rob.scala 147:39]
  wire  _GEN_27847 = io_i_ex_res_packs_1_valid ? _GEN_25671 : _GEN_23495; // @[rob.scala 147:39]
  wire  _GEN_27848 = io_i_ex_res_packs_1_valid ? _GEN_25672 : _GEN_23496; // @[rob.scala 147:39]
  wire  _GEN_27849 = io_i_ex_res_packs_1_valid ? _GEN_25673 : _GEN_23497; // @[rob.scala 147:39]
  wire  _GEN_27850 = io_i_ex_res_packs_1_valid ? _GEN_25674 : _GEN_23498; // @[rob.scala 147:39]
  wire  _GEN_27851 = io_i_ex_res_packs_1_valid ? _GEN_25675 : _GEN_23499; // @[rob.scala 147:39]
  wire  _GEN_27852 = io_i_ex_res_packs_1_valid ? _GEN_25676 : _GEN_23500; // @[rob.scala 147:39]
  wire  _GEN_27853 = io_i_ex_res_packs_1_valid ? _GEN_25677 : _GEN_23501; // @[rob.scala 147:39]
  wire  _GEN_27854 = io_i_ex_res_packs_1_valid ? _GEN_25678 : _GEN_23502; // @[rob.scala 147:39]
  wire  _GEN_27855 = io_i_ex_res_packs_1_valid ? _GEN_25679 : _GEN_23503; // @[rob.scala 147:39]
  wire  _GEN_27856 = io_i_ex_res_packs_1_valid ? _GEN_25680 : _GEN_23504; // @[rob.scala 147:39]
  wire  _GEN_27857 = io_i_ex_res_packs_1_valid ? _GEN_25681 : _GEN_23505; // @[rob.scala 147:39]
  wire  _GEN_27858 = io_i_ex_res_packs_1_valid ? _GEN_25682 : _GEN_23506; // @[rob.scala 147:39]
  wire  _GEN_27859 = io_i_ex_res_packs_1_valid ? _GEN_25683 : _GEN_23507; // @[rob.scala 147:39]
  wire  _GEN_27860 = io_i_ex_res_packs_1_valid ? _GEN_25684 : _GEN_23508; // @[rob.scala 147:39]
  wire  _GEN_27861 = io_i_ex_res_packs_1_valid ? _GEN_25685 : _GEN_23509; // @[rob.scala 147:39]
  wire  _GEN_27862 = io_i_ex_res_packs_1_valid ? _GEN_25686 : _GEN_23510; // @[rob.scala 147:39]
  wire  _GEN_27863 = io_i_ex_res_packs_1_valid ? _GEN_25687 : _GEN_23511; // @[rob.scala 147:39]
  wire  _GEN_27864 = io_i_ex_res_packs_1_valid ? _GEN_25688 : _GEN_23512; // @[rob.scala 147:39]
  wire  _GEN_27865 = io_i_ex_res_packs_1_valid ? _GEN_25689 : _GEN_23513; // @[rob.scala 147:39]
  wire  _GEN_27866 = io_i_ex_res_packs_1_valid ? _GEN_25690 : _GEN_23514; // @[rob.scala 147:39]
  wire  _GEN_27867 = io_i_ex_res_packs_1_valid ? _GEN_25691 : _GEN_23515; // @[rob.scala 147:39]
  wire  _GEN_27868 = io_i_ex_res_packs_1_valid ? _GEN_25692 : _GEN_23516; // @[rob.scala 147:39]
  wire  _GEN_27869 = io_i_ex_res_packs_1_valid ? _GEN_25693 : _GEN_23517; // @[rob.scala 147:39]
  wire  _GEN_27870 = io_i_ex_res_packs_1_valid ? _GEN_25694 : _GEN_23518; // @[rob.scala 147:39]
  wire  _GEN_27871 = io_i_ex_res_packs_1_valid ? _GEN_25695 : _GEN_23519; // @[rob.scala 147:39]
  wire  _GEN_27872 = io_i_ex_res_packs_1_valid ? _GEN_25696 : _GEN_23520; // @[rob.scala 147:39]
  wire  _GEN_27873 = io_i_ex_res_packs_1_valid ? _GEN_25697 : _GEN_23521; // @[rob.scala 147:39]
  wire  _GEN_27874 = io_i_ex_res_packs_1_valid ? _GEN_25698 : _GEN_23522; // @[rob.scala 147:39]
  wire  _GEN_27875 = io_i_ex_res_packs_1_valid ? _GEN_25699 : _GEN_23523; // @[rob.scala 147:39]
  wire  _GEN_27876 = io_i_ex_res_packs_1_valid ? _GEN_25700 : _GEN_23524; // @[rob.scala 147:39]
  wire  _GEN_27877 = io_i_ex_res_packs_1_valid ? _GEN_25701 : _GEN_23525; // @[rob.scala 147:39]
  wire  _GEN_27878 = io_i_ex_res_packs_1_valid ? _GEN_25702 : _GEN_23526; // @[rob.scala 147:39]
  wire  _GEN_27879 = io_i_ex_res_packs_1_valid ? _GEN_25703 : _GEN_23527; // @[rob.scala 147:39]
  wire  _GEN_27880 = io_i_ex_res_packs_1_valid ? _GEN_25704 : _GEN_23528; // @[rob.scala 147:39]
  wire  _GEN_27881 = io_i_ex_res_packs_1_valid ? _GEN_25705 : _GEN_23529; // @[rob.scala 147:39]
  wire  _GEN_27882 = io_i_ex_res_packs_1_valid ? _GEN_25706 : _GEN_23530; // @[rob.scala 147:39]
  wire  _GEN_27883 = io_i_ex_res_packs_1_valid ? _GEN_25707 : _GEN_23531; // @[rob.scala 147:39]
  wire  _GEN_27884 = io_i_ex_res_packs_1_valid ? _GEN_25708 : _GEN_23532; // @[rob.scala 147:39]
  wire  _GEN_27885 = io_i_ex_res_packs_1_valid ? _GEN_25709 : _GEN_23533; // @[rob.scala 147:39]
  wire  _GEN_27886 = io_i_ex_res_packs_1_valid ? _GEN_25710 : _GEN_23534; // @[rob.scala 147:39]
  wire  _GEN_27887 = io_i_ex_res_packs_1_valid ? _GEN_25711 : _GEN_23535; // @[rob.scala 147:39]
  wire  _GEN_27888 = io_i_ex_res_packs_1_valid ? _GEN_25712 : _GEN_23536; // @[rob.scala 147:39]
  wire  _GEN_27889 = io_i_ex_res_packs_1_valid ? _GEN_25713 : _GEN_23537; // @[rob.scala 147:39]
  wire  _GEN_27890 = io_i_ex_res_packs_1_valid ? _GEN_25714 : _GEN_23538; // @[rob.scala 147:39]
  wire  _GEN_27891 = io_i_ex_res_packs_1_valid ? _GEN_25715 : _GEN_23539; // @[rob.scala 147:39]
  wire  _GEN_27892 = io_i_ex_res_packs_1_valid ? _GEN_25716 : _GEN_23540; // @[rob.scala 147:39]
  wire  _GEN_27893 = io_i_ex_res_packs_1_valid ? _GEN_25717 : _GEN_23541; // @[rob.scala 147:39]
  wire  _GEN_27894 = io_i_ex_res_packs_1_valid ? _GEN_25718 : _GEN_23542; // @[rob.scala 147:39]
  wire  _GEN_27895 = io_i_ex_res_packs_1_valid ? _GEN_25719 : _GEN_23543; // @[rob.scala 147:39]
  wire  _GEN_27896 = io_i_ex_res_packs_1_valid ? _GEN_25720 : _GEN_23544; // @[rob.scala 147:39]
  wire  _GEN_27897 = io_i_ex_res_packs_1_valid ? _GEN_25721 : _GEN_23545; // @[rob.scala 147:39]
  wire  _GEN_27898 = io_i_ex_res_packs_1_valid ? _GEN_25722 : _GEN_23546; // @[rob.scala 147:39]
  wire  _GEN_27899 = io_i_ex_res_packs_1_valid ? _GEN_25723 : _GEN_23547; // @[rob.scala 147:39]
  wire  _GEN_27900 = io_i_ex_res_packs_1_valid ? _GEN_25724 : _GEN_23548; // @[rob.scala 147:39]
  wire  _GEN_27901 = io_i_ex_res_packs_1_valid ? _GEN_25725 : _GEN_23549; // @[rob.scala 147:39]
  wire  _GEN_27902 = io_i_ex_res_packs_1_valid ? _GEN_25726 : _GEN_23550; // @[rob.scala 147:39]
  wire  _GEN_27903 = io_i_ex_res_packs_1_valid ? _GEN_25727 : _GEN_23551; // @[rob.scala 147:39]
  wire  _GEN_27904 = io_i_ex_res_packs_1_valid ? _GEN_25728 : _GEN_23552; // @[rob.scala 147:39]
  wire  _GEN_27905 = io_i_ex_res_packs_1_valid ? _GEN_25729 : _GEN_23553; // @[rob.scala 147:39]
  wire  _T_26 = next_will_commit_0 & next_will_commit_1; // @[rob.scala 155:32]
  wire  _GEN_27906 = 6'h0 == commit_ptr[5:0] ? 1'h0 : _GEN_25730; // @[rob.scala 156:{31,31}]
  wire  _GEN_27907 = 6'h1 == commit_ptr[5:0] ? 1'h0 : _GEN_25731; // @[rob.scala 156:{31,31}]
  wire  _GEN_27908 = 6'h2 == commit_ptr[5:0] ? 1'h0 : _GEN_25732; // @[rob.scala 156:{31,31}]
  wire  _GEN_27909 = 6'h3 == commit_ptr[5:0] ? 1'h0 : _GEN_25733; // @[rob.scala 156:{31,31}]
  wire  _GEN_27910 = 6'h4 == commit_ptr[5:0] ? 1'h0 : _GEN_25734; // @[rob.scala 156:{31,31}]
  wire  _GEN_27911 = 6'h5 == commit_ptr[5:0] ? 1'h0 : _GEN_25735; // @[rob.scala 156:{31,31}]
  wire  _GEN_27912 = 6'h6 == commit_ptr[5:0] ? 1'h0 : _GEN_25736; // @[rob.scala 156:{31,31}]
  wire  _GEN_27913 = 6'h7 == commit_ptr[5:0] ? 1'h0 : _GEN_25737; // @[rob.scala 156:{31,31}]
  wire  _GEN_27914 = 6'h8 == commit_ptr[5:0] ? 1'h0 : _GEN_25738; // @[rob.scala 156:{31,31}]
  wire  _GEN_27915 = 6'h9 == commit_ptr[5:0] ? 1'h0 : _GEN_25739; // @[rob.scala 156:{31,31}]
  wire  _GEN_27916 = 6'ha == commit_ptr[5:0] ? 1'h0 : _GEN_25740; // @[rob.scala 156:{31,31}]
  wire  _GEN_27917 = 6'hb == commit_ptr[5:0] ? 1'h0 : _GEN_25741; // @[rob.scala 156:{31,31}]
  wire  _GEN_27918 = 6'hc == commit_ptr[5:0] ? 1'h0 : _GEN_25742; // @[rob.scala 156:{31,31}]
  wire  _GEN_27919 = 6'hd == commit_ptr[5:0] ? 1'h0 : _GEN_25743; // @[rob.scala 156:{31,31}]
  wire  _GEN_27920 = 6'he == commit_ptr[5:0] ? 1'h0 : _GEN_25744; // @[rob.scala 156:{31,31}]
  wire  _GEN_27921 = 6'hf == commit_ptr[5:0] ? 1'h0 : _GEN_25745; // @[rob.scala 156:{31,31}]
  wire  _GEN_27922 = 6'h10 == commit_ptr[5:0] ? 1'h0 : _GEN_25746; // @[rob.scala 156:{31,31}]
  wire  _GEN_27923 = 6'h11 == commit_ptr[5:0] ? 1'h0 : _GEN_25747; // @[rob.scala 156:{31,31}]
  wire  _GEN_27924 = 6'h12 == commit_ptr[5:0] ? 1'h0 : _GEN_25748; // @[rob.scala 156:{31,31}]
  wire  _GEN_27925 = 6'h13 == commit_ptr[5:0] ? 1'h0 : _GEN_25749; // @[rob.scala 156:{31,31}]
  wire  _GEN_27926 = 6'h14 == commit_ptr[5:0] ? 1'h0 : _GEN_25750; // @[rob.scala 156:{31,31}]
  wire  _GEN_27927 = 6'h15 == commit_ptr[5:0] ? 1'h0 : _GEN_25751; // @[rob.scala 156:{31,31}]
  wire  _GEN_27928 = 6'h16 == commit_ptr[5:0] ? 1'h0 : _GEN_25752; // @[rob.scala 156:{31,31}]
  wire  _GEN_27929 = 6'h17 == commit_ptr[5:0] ? 1'h0 : _GEN_25753; // @[rob.scala 156:{31,31}]
  wire  _GEN_27930 = 6'h18 == commit_ptr[5:0] ? 1'h0 : _GEN_25754; // @[rob.scala 156:{31,31}]
  wire  _GEN_27931 = 6'h19 == commit_ptr[5:0] ? 1'h0 : _GEN_25755; // @[rob.scala 156:{31,31}]
  wire  _GEN_27932 = 6'h1a == commit_ptr[5:0] ? 1'h0 : _GEN_25756; // @[rob.scala 156:{31,31}]
  wire  _GEN_27933 = 6'h1b == commit_ptr[5:0] ? 1'h0 : _GEN_25757; // @[rob.scala 156:{31,31}]
  wire  _GEN_27934 = 6'h1c == commit_ptr[5:0] ? 1'h0 : _GEN_25758; // @[rob.scala 156:{31,31}]
  wire  _GEN_27935 = 6'h1d == commit_ptr[5:0] ? 1'h0 : _GEN_25759; // @[rob.scala 156:{31,31}]
  wire  _GEN_27936 = 6'h1e == commit_ptr[5:0] ? 1'h0 : _GEN_25760; // @[rob.scala 156:{31,31}]
  wire  _GEN_27937 = 6'h1f == commit_ptr[5:0] ? 1'h0 : _GEN_25761; // @[rob.scala 156:{31,31}]
  wire  _GEN_27938 = 6'h20 == commit_ptr[5:0] ? 1'h0 : _GEN_25762; // @[rob.scala 156:{31,31}]
  wire  _GEN_27939 = 6'h21 == commit_ptr[5:0] ? 1'h0 : _GEN_25763; // @[rob.scala 156:{31,31}]
  wire  _GEN_27940 = 6'h22 == commit_ptr[5:0] ? 1'h0 : _GEN_25764; // @[rob.scala 156:{31,31}]
  wire  _GEN_27941 = 6'h23 == commit_ptr[5:0] ? 1'h0 : _GEN_25765; // @[rob.scala 156:{31,31}]
  wire  _GEN_27942 = 6'h24 == commit_ptr[5:0] ? 1'h0 : _GEN_25766; // @[rob.scala 156:{31,31}]
  wire  _GEN_27943 = 6'h25 == commit_ptr[5:0] ? 1'h0 : _GEN_25767; // @[rob.scala 156:{31,31}]
  wire  _GEN_27944 = 6'h26 == commit_ptr[5:0] ? 1'h0 : _GEN_25768; // @[rob.scala 156:{31,31}]
  wire  _GEN_27945 = 6'h27 == commit_ptr[5:0] ? 1'h0 : _GEN_25769; // @[rob.scala 156:{31,31}]
  wire  _GEN_27946 = 6'h28 == commit_ptr[5:0] ? 1'h0 : _GEN_25770; // @[rob.scala 156:{31,31}]
  wire  _GEN_27947 = 6'h29 == commit_ptr[5:0] ? 1'h0 : _GEN_25771; // @[rob.scala 156:{31,31}]
  wire  _GEN_27948 = 6'h2a == commit_ptr[5:0] ? 1'h0 : _GEN_25772; // @[rob.scala 156:{31,31}]
  wire  _GEN_27949 = 6'h2b == commit_ptr[5:0] ? 1'h0 : _GEN_25773; // @[rob.scala 156:{31,31}]
  wire  _GEN_27950 = 6'h2c == commit_ptr[5:0] ? 1'h0 : _GEN_25774; // @[rob.scala 156:{31,31}]
  wire  _GEN_27951 = 6'h2d == commit_ptr[5:0] ? 1'h0 : _GEN_25775; // @[rob.scala 156:{31,31}]
  wire  _GEN_27952 = 6'h2e == commit_ptr[5:0] ? 1'h0 : _GEN_25776; // @[rob.scala 156:{31,31}]
  wire  _GEN_27953 = 6'h2f == commit_ptr[5:0] ? 1'h0 : _GEN_25777; // @[rob.scala 156:{31,31}]
  wire  _GEN_27954 = 6'h30 == commit_ptr[5:0] ? 1'h0 : _GEN_25778; // @[rob.scala 156:{31,31}]
  wire  _GEN_27955 = 6'h31 == commit_ptr[5:0] ? 1'h0 : _GEN_25779; // @[rob.scala 156:{31,31}]
  wire  _GEN_27956 = 6'h32 == commit_ptr[5:0] ? 1'h0 : _GEN_25780; // @[rob.scala 156:{31,31}]
  wire  _GEN_27957 = 6'h33 == commit_ptr[5:0] ? 1'h0 : _GEN_25781; // @[rob.scala 156:{31,31}]
  wire  _GEN_27958 = 6'h34 == commit_ptr[5:0] ? 1'h0 : _GEN_25782; // @[rob.scala 156:{31,31}]
  wire  _GEN_27959 = 6'h35 == commit_ptr[5:0] ? 1'h0 : _GEN_25783; // @[rob.scala 156:{31,31}]
  wire  _GEN_27960 = 6'h36 == commit_ptr[5:0] ? 1'h0 : _GEN_25784; // @[rob.scala 156:{31,31}]
  wire  _GEN_27961 = 6'h37 == commit_ptr[5:0] ? 1'h0 : _GEN_25785; // @[rob.scala 156:{31,31}]
  wire  _GEN_27962 = 6'h38 == commit_ptr[5:0] ? 1'h0 : _GEN_25786; // @[rob.scala 156:{31,31}]
  wire  _GEN_27963 = 6'h39 == commit_ptr[5:0] ? 1'h0 : _GEN_25787; // @[rob.scala 156:{31,31}]
  wire  _GEN_27964 = 6'h3a == commit_ptr[5:0] ? 1'h0 : _GEN_25788; // @[rob.scala 156:{31,31}]
  wire  _GEN_27965 = 6'h3b == commit_ptr[5:0] ? 1'h0 : _GEN_25789; // @[rob.scala 156:{31,31}]
  wire  _GEN_27966 = 6'h3c == commit_ptr[5:0] ? 1'h0 : _GEN_25790; // @[rob.scala 156:{31,31}]
  wire  _GEN_27967 = 6'h3d == commit_ptr[5:0] ? 1'h0 : _GEN_25791; // @[rob.scala 156:{31,31}]
  wire  _GEN_27968 = 6'h3e == commit_ptr[5:0] ? 1'h0 : _GEN_25792; // @[rob.scala 156:{31,31}]
  wire  _GEN_27969 = 6'h3f == commit_ptr[5:0] ? 1'h0 : _GEN_25793; // @[rob.scala 156:{31,31}]
  wire  _GEN_27970 = 6'h0 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27906; // @[rob.scala 157:{35,35}]
  wire  _GEN_27971 = 6'h1 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27907; // @[rob.scala 157:{35,35}]
  wire  _GEN_27972 = 6'h2 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27908; // @[rob.scala 157:{35,35}]
  wire  _GEN_27973 = 6'h3 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27909; // @[rob.scala 157:{35,35}]
  wire  _GEN_27974 = 6'h4 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27910; // @[rob.scala 157:{35,35}]
  wire  _GEN_27975 = 6'h5 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27911; // @[rob.scala 157:{35,35}]
  wire  _GEN_27976 = 6'h6 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27912; // @[rob.scala 157:{35,35}]
  wire  _GEN_27977 = 6'h7 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27913; // @[rob.scala 157:{35,35}]
  wire  _GEN_27978 = 6'h8 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27914; // @[rob.scala 157:{35,35}]
  wire  _GEN_27979 = 6'h9 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27915; // @[rob.scala 157:{35,35}]
  wire  _GEN_27980 = 6'ha == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27916; // @[rob.scala 157:{35,35}]
  wire  _GEN_27981 = 6'hb == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27917; // @[rob.scala 157:{35,35}]
  wire  _GEN_27982 = 6'hc == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27918; // @[rob.scala 157:{35,35}]
  wire  _GEN_27983 = 6'hd == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27919; // @[rob.scala 157:{35,35}]
  wire  _GEN_27984 = 6'he == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27920; // @[rob.scala 157:{35,35}]
  wire  _GEN_27985 = 6'hf == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27921; // @[rob.scala 157:{35,35}]
  wire  _GEN_27986 = 6'h10 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27922; // @[rob.scala 157:{35,35}]
  wire  _GEN_27987 = 6'h11 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27923; // @[rob.scala 157:{35,35}]
  wire  _GEN_27988 = 6'h12 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27924; // @[rob.scala 157:{35,35}]
  wire  _GEN_27989 = 6'h13 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27925; // @[rob.scala 157:{35,35}]
  wire  _GEN_27990 = 6'h14 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27926; // @[rob.scala 157:{35,35}]
  wire  _GEN_27991 = 6'h15 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27927; // @[rob.scala 157:{35,35}]
  wire  _GEN_27992 = 6'h16 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27928; // @[rob.scala 157:{35,35}]
  wire  _GEN_27993 = 6'h17 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27929; // @[rob.scala 157:{35,35}]
  wire  _GEN_27994 = 6'h18 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27930; // @[rob.scala 157:{35,35}]
  wire  _GEN_27995 = 6'h19 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27931; // @[rob.scala 157:{35,35}]
  wire  _GEN_27996 = 6'h1a == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27932; // @[rob.scala 157:{35,35}]
  wire  _GEN_27997 = 6'h1b == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27933; // @[rob.scala 157:{35,35}]
  wire  _GEN_27998 = 6'h1c == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27934; // @[rob.scala 157:{35,35}]
  wire  _GEN_27999 = 6'h1d == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27935; // @[rob.scala 157:{35,35}]
  wire  _GEN_28000 = 6'h1e == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27936; // @[rob.scala 157:{35,35}]
  wire  _GEN_28001 = 6'h1f == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27937; // @[rob.scala 157:{35,35}]
  wire  _GEN_28002 = 6'h20 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27938; // @[rob.scala 157:{35,35}]
  wire  _GEN_28003 = 6'h21 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27939; // @[rob.scala 157:{35,35}]
  wire  _GEN_28004 = 6'h22 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27940; // @[rob.scala 157:{35,35}]
  wire  _GEN_28005 = 6'h23 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27941; // @[rob.scala 157:{35,35}]
  wire  _GEN_28006 = 6'h24 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27942; // @[rob.scala 157:{35,35}]
  wire  _GEN_28007 = 6'h25 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27943; // @[rob.scala 157:{35,35}]
  wire  _GEN_28008 = 6'h26 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27944; // @[rob.scala 157:{35,35}]
  wire  _GEN_28009 = 6'h27 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27945; // @[rob.scala 157:{35,35}]
  wire  _GEN_28010 = 6'h28 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27946; // @[rob.scala 157:{35,35}]
  wire  _GEN_28011 = 6'h29 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27947; // @[rob.scala 157:{35,35}]
  wire  _GEN_28012 = 6'h2a == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27948; // @[rob.scala 157:{35,35}]
  wire  _GEN_28013 = 6'h2b == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27949; // @[rob.scala 157:{35,35}]
  wire  _GEN_28014 = 6'h2c == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27950; // @[rob.scala 157:{35,35}]
  wire  _GEN_28015 = 6'h2d == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27951; // @[rob.scala 157:{35,35}]
  wire  _GEN_28016 = 6'h2e == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27952; // @[rob.scala 157:{35,35}]
  wire  _GEN_28017 = 6'h2f == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27953; // @[rob.scala 157:{35,35}]
  wire  _GEN_28018 = 6'h30 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27954; // @[rob.scala 157:{35,35}]
  wire  _GEN_28019 = 6'h31 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27955; // @[rob.scala 157:{35,35}]
  wire  _GEN_28020 = 6'h32 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27956; // @[rob.scala 157:{35,35}]
  wire  _GEN_28021 = 6'h33 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27957; // @[rob.scala 157:{35,35}]
  wire  _GEN_28022 = 6'h34 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27958; // @[rob.scala 157:{35,35}]
  wire  _GEN_28023 = 6'h35 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27959; // @[rob.scala 157:{35,35}]
  wire  _GEN_28024 = 6'h36 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27960; // @[rob.scala 157:{35,35}]
  wire  _GEN_28025 = 6'h37 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27961; // @[rob.scala 157:{35,35}]
  wire  _GEN_28026 = 6'h38 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27962; // @[rob.scala 157:{35,35}]
  wire  _GEN_28027 = 6'h39 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27963; // @[rob.scala 157:{35,35}]
  wire  _GEN_28028 = 6'h3a == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27964; // @[rob.scala 157:{35,35}]
  wire  _GEN_28029 = 6'h3b == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27965; // @[rob.scala 157:{35,35}]
  wire  _GEN_28030 = 6'h3c == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27966; // @[rob.scala 157:{35,35}]
  wire  _GEN_28031 = 6'h3d == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27967; // @[rob.scala 157:{35,35}]
  wire  _GEN_28032 = 6'h3e == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27968; // @[rob.scala 157:{35,35}]
  wire  _GEN_28033 = 6'h3f == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_27969; // @[rob.scala 157:{35,35}]
  wire [6:0] _commit_ptr_T_1 = commit_ptr + 7'h2; // @[rob.scala 158:34]
  wire  _GEN_28098 = next_will_commit_0 ? _GEN_27906 : _GEN_25730; // @[rob.scala 159:38]
  wire  _GEN_28099 = next_will_commit_0 ? _GEN_27907 : _GEN_25731; // @[rob.scala 159:38]
  wire  _GEN_28100 = next_will_commit_0 ? _GEN_27908 : _GEN_25732; // @[rob.scala 159:38]
  wire  _GEN_28101 = next_will_commit_0 ? _GEN_27909 : _GEN_25733; // @[rob.scala 159:38]
  wire  _GEN_28102 = next_will_commit_0 ? _GEN_27910 : _GEN_25734; // @[rob.scala 159:38]
  wire  _GEN_28103 = next_will_commit_0 ? _GEN_27911 : _GEN_25735; // @[rob.scala 159:38]
  wire  _GEN_28104 = next_will_commit_0 ? _GEN_27912 : _GEN_25736; // @[rob.scala 159:38]
  wire  _GEN_28105 = next_will_commit_0 ? _GEN_27913 : _GEN_25737; // @[rob.scala 159:38]
  wire  _GEN_28106 = next_will_commit_0 ? _GEN_27914 : _GEN_25738; // @[rob.scala 159:38]
  wire  _GEN_28107 = next_will_commit_0 ? _GEN_27915 : _GEN_25739; // @[rob.scala 159:38]
  wire  _GEN_28108 = next_will_commit_0 ? _GEN_27916 : _GEN_25740; // @[rob.scala 159:38]
  wire  _GEN_28109 = next_will_commit_0 ? _GEN_27917 : _GEN_25741; // @[rob.scala 159:38]
  wire  _GEN_28110 = next_will_commit_0 ? _GEN_27918 : _GEN_25742; // @[rob.scala 159:38]
  wire  _GEN_28111 = next_will_commit_0 ? _GEN_27919 : _GEN_25743; // @[rob.scala 159:38]
  wire  _GEN_28112 = next_will_commit_0 ? _GEN_27920 : _GEN_25744; // @[rob.scala 159:38]
  wire  _GEN_28113 = next_will_commit_0 ? _GEN_27921 : _GEN_25745; // @[rob.scala 159:38]
  wire  _GEN_28114 = next_will_commit_0 ? _GEN_27922 : _GEN_25746; // @[rob.scala 159:38]
  wire  _GEN_28115 = next_will_commit_0 ? _GEN_27923 : _GEN_25747; // @[rob.scala 159:38]
  wire  _GEN_28116 = next_will_commit_0 ? _GEN_27924 : _GEN_25748; // @[rob.scala 159:38]
  wire  _GEN_28117 = next_will_commit_0 ? _GEN_27925 : _GEN_25749; // @[rob.scala 159:38]
  wire  _GEN_28118 = next_will_commit_0 ? _GEN_27926 : _GEN_25750; // @[rob.scala 159:38]
  wire  _GEN_28119 = next_will_commit_0 ? _GEN_27927 : _GEN_25751; // @[rob.scala 159:38]
  wire  _GEN_28120 = next_will_commit_0 ? _GEN_27928 : _GEN_25752; // @[rob.scala 159:38]
  wire  _GEN_28121 = next_will_commit_0 ? _GEN_27929 : _GEN_25753; // @[rob.scala 159:38]
  wire  _GEN_28122 = next_will_commit_0 ? _GEN_27930 : _GEN_25754; // @[rob.scala 159:38]
  wire  _GEN_28123 = next_will_commit_0 ? _GEN_27931 : _GEN_25755; // @[rob.scala 159:38]
  wire  _GEN_28124 = next_will_commit_0 ? _GEN_27932 : _GEN_25756; // @[rob.scala 159:38]
  wire  _GEN_28125 = next_will_commit_0 ? _GEN_27933 : _GEN_25757; // @[rob.scala 159:38]
  wire  _GEN_28126 = next_will_commit_0 ? _GEN_27934 : _GEN_25758; // @[rob.scala 159:38]
  wire  _GEN_28127 = next_will_commit_0 ? _GEN_27935 : _GEN_25759; // @[rob.scala 159:38]
  wire  _GEN_28128 = next_will_commit_0 ? _GEN_27936 : _GEN_25760; // @[rob.scala 159:38]
  wire  _GEN_28129 = next_will_commit_0 ? _GEN_27937 : _GEN_25761; // @[rob.scala 159:38]
  wire  _GEN_28130 = next_will_commit_0 ? _GEN_27938 : _GEN_25762; // @[rob.scala 159:38]
  wire  _GEN_28131 = next_will_commit_0 ? _GEN_27939 : _GEN_25763; // @[rob.scala 159:38]
  wire  _GEN_28132 = next_will_commit_0 ? _GEN_27940 : _GEN_25764; // @[rob.scala 159:38]
  wire  _GEN_28133 = next_will_commit_0 ? _GEN_27941 : _GEN_25765; // @[rob.scala 159:38]
  wire  _GEN_28134 = next_will_commit_0 ? _GEN_27942 : _GEN_25766; // @[rob.scala 159:38]
  wire  _GEN_28135 = next_will_commit_0 ? _GEN_27943 : _GEN_25767; // @[rob.scala 159:38]
  wire  _GEN_28136 = next_will_commit_0 ? _GEN_27944 : _GEN_25768; // @[rob.scala 159:38]
  wire  _GEN_28137 = next_will_commit_0 ? _GEN_27945 : _GEN_25769; // @[rob.scala 159:38]
  wire  _GEN_28138 = next_will_commit_0 ? _GEN_27946 : _GEN_25770; // @[rob.scala 159:38]
  wire  _GEN_28139 = next_will_commit_0 ? _GEN_27947 : _GEN_25771; // @[rob.scala 159:38]
  wire  _GEN_28140 = next_will_commit_0 ? _GEN_27948 : _GEN_25772; // @[rob.scala 159:38]
  wire  _GEN_28141 = next_will_commit_0 ? _GEN_27949 : _GEN_25773; // @[rob.scala 159:38]
  wire  _GEN_28142 = next_will_commit_0 ? _GEN_27950 : _GEN_25774; // @[rob.scala 159:38]
  wire  _GEN_28143 = next_will_commit_0 ? _GEN_27951 : _GEN_25775; // @[rob.scala 159:38]
  wire  _GEN_28144 = next_will_commit_0 ? _GEN_27952 : _GEN_25776; // @[rob.scala 159:38]
  wire  _GEN_28145 = next_will_commit_0 ? _GEN_27953 : _GEN_25777; // @[rob.scala 159:38]
  wire  _GEN_28146 = next_will_commit_0 ? _GEN_27954 : _GEN_25778; // @[rob.scala 159:38]
  wire  _GEN_28147 = next_will_commit_0 ? _GEN_27955 : _GEN_25779; // @[rob.scala 159:38]
  wire  _GEN_28148 = next_will_commit_0 ? _GEN_27956 : _GEN_25780; // @[rob.scala 159:38]
  wire  _GEN_28149 = next_will_commit_0 ? _GEN_27957 : _GEN_25781; // @[rob.scala 159:38]
  wire  _GEN_28150 = next_will_commit_0 ? _GEN_27958 : _GEN_25782; // @[rob.scala 159:38]
  wire  _GEN_28151 = next_will_commit_0 ? _GEN_27959 : _GEN_25783; // @[rob.scala 159:38]
  wire  _GEN_28152 = next_will_commit_0 ? _GEN_27960 : _GEN_25784; // @[rob.scala 159:38]
  wire  _GEN_28153 = next_will_commit_0 ? _GEN_27961 : _GEN_25785; // @[rob.scala 159:38]
  wire  _GEN_28154 = next_will_commit_0 ? _GEN_27962 : _GEN_25786; // @[rob.scala 159:38]
  wire  _GEN_28155 = next_will_commit_0 ? _GEN_27963 : _GEN_25787; // @[rob.scala 159:38]
  wire  _GEN_28156 = next_will_commit_0 ? _GEN_27964 : _GEN_25788; // @[rob.scala 159:38]
  wire  _GEN_28157 = next_will_commit_0 ? _GEN_27965 : _GEN_25789; // @[rob.scala 159:38]
  wire  _GEN_28158 = next_will_commit_0 ? _GEN_27966 : _GEN_25790; // @[rob.scala 159:38]
  wire  _GEN_28159 = next_will_commit_0 ? _GEN_27967 : _GEN_25791; // @[rob.scala 159:38]
  wire  _GEN_28160 = next_will_commit_0 ? _GEN_27968 : _GEN_25792; // @[rob.scala 159:38]
  wire  _GEN_28161 = next_will_commit_0 ? _GEN_27969 : _GEN_25793; // @[rob.scala 159:38]
  wire [6:0] _GEN_28162 = next_will_commit_0 ? _next_can_commit_1_T_1 : commit_ptr; // @[rob.scala 159:38 161:20 46:29]
  wire  _GEN_28163 = next_will_commit_0 & next_will_commit_1 ? _GEN_27970 : _GEN_28098; // @[rob.scala 155:55]
  wire  _GEN_28164 = next_will_commit_0 & next_will_commit_1 ? _GEN_27971 : _GEN_28099; // @[rob.scala 155:55]
  wire  _GEN_28165 = next_will_commit_0 & next_will_commit_1 ? _GEN_27972 : _GEN_28100; // @[rob.scala 155:55]
  wire  _GEN_28166 = next_will_commit_0 & next_will_commit_1 ? _GEN_27973 : _GEN_28101; // @[rob.scala 155:55]
  wire  _GEN_28167 = next_will_commit_0 & next_will_commit_1 ? _GEN_27974 : _GEN_28102; // @[rob.scala 155:55]
  wire  _GEN_28168 = next_will_commit_0 & next_will_commit_1 ? _GEN_27975 : _GEN_28103; // @[rob.scala 155:55]
  wire  _GEN_28169 = next_will_commit_0 & next_will_commit_1 ? _GEN_27976 : _GEN_28104; // @[rob.scala 155:55]
  wire  _GEN_28170 = next_will_commit_0 & next_will_commit_1 ? _GEN_27977 : _GEN_28105; // @[rob.scala 155:55]
  wire  _GEN_28171 = next_will_commit_0 & next_will_commit_1 ? _GEN_27978 : _GEN_28106; // @[rob.scala 155:55]
  wire  _GEN_28172 = next_will_commit_0 & next_will_commit_1 ? _GEN_27979 : _GEN_28107; // @[rob.scala 155:55]
  wire  _GEN_28173 = next_will_commit_0 & next_will_commit_1 ? _GEN_27980 : _GEN_28108; // @[rob.scala 155:55]
  wire  _GEN_28174 = next_will_commit_0 & next_will_commit_1 ? _GEN_27981 : _GEN_28109; // @[rob.scala 155:55]
  wire  _GEN_28175 = next_will_commit_0 & next_will_commit_1 ? _GEN_27982 : _GEN_28110; // @[rob.scala 155:55]
  wire  _GEN_28176 = next_will_commit_0 & next_will_commit_1 ? _GEN_27983 : _GEN_28111; // @[rob.scala 155:55]
  wire  _GEN_28177 = next_will_commit_0 & next_will_commit_1 ? _GEN_27984 : _GEN_28112; // @[rob.scala 155:55]
  wire  _GEN_28178 = next_will_commit_0 & next_will_commit_1 ? _GEN_27985 : _GEN_28113; // @[rob.scala 155:55]
  wire  _GEN_28179 = next_will_commit_0 & next_will_commit_1 ? _GEN_27986 : _GEN_28114; // @[rob.scala 155:55]
  wire  _GEN_28180 = next_will_commit_0 & next_will_commit_1 ? _GEN_27987 : _GEN_28115; // @[rob.scala 155:55]
  wire  _GEN_28181 = next_will_commit_0 & next_will_commit_1 ? _GEN_27988 : _GEN_28116; // @[rob.scala 155:55]
  wire  _GEN_28182 = next_will_commit_0 & next_will_commit_1 ? _GEN_27989 : _GEN_28117; // @[rob.scala 155:55]
  wire  _GEN_28183 = next_will_commit_0 & next_will_commit_1 ? _GEN_27990 : _GEN_28118; // @[rob.scala 155:55]
  wire  _GEN_28184 = next_will_commit_0 & next_will_commit_1 ? _GEN_27991 : _GEN_28119; // @[rob.scala 155:55]
  wire  _GEN_28185 = next_will_commit_0 & next_will_commit_1 ? _GEN_27992 : _GEN_28120; // @[rob.scala 155:55]
  wire  _GEN_28186 = next_will_commit_0 & next_will_commit_1 ? _GEN_27993 : _GEN_28121; // @[rob.scala 155:55]
  wire  _GEN_28187 = next_will_commit_0 & next_will_commit_1 ? _GEN_27994 : _GEN_28122; // @[rob.scala 155:55]
  wire  _GEN_28188 = next_will_commit_0 & next_will_commit_1 ? _GEN_27995 : _GEN_28123; // @[rob.scala 155:55]
  wire  _GEN_28189 = next_will_commit_0 & next_will_commit_1 ? _GEN_27996 : _GEN_28124; // @[rob.scala 155:55]
  wire  _GEN_28190 = next_will_commit_0 & next_will_commit_1 ? _GEN_27997 : _GEN_28125; // @[rob.scala 155:55]
  wire  _GEN_28191 = next_will_commit_0 & next_will_commit_1 ? _GEN_27998 : _GEN_28126; // @[rob.scala 155:55]
  wire  _GEN_28192 = next_will_commit_0 & next_will_commit_1 ? _GEN_27999 : _GEN_28127; // @[rob.scala 155:55]
  wire  _GEN_28193 = next_will_commit_0 & next_will_commit_1 ? _GEN_28000 : _GEN_28128; // @[rob.scala 155:55]
  wire  _GEN_28194 = next_will_commit_0 & next_will_commit_1 ? _GEN_28001 : _GEN_28129; // @[rob.scala 155:55]
  wire  _GEN_28195 = next_will_commit_0 & next_will_commit_1 ? _GEN_28002 : _GEN_28130; // @[rob.scala 155:55]
  wire  _GEN_28196 = next_will_commit_0 & next_will_commit_1 ? _GEN_28003 : _GEN_28131; // @[rob.scala 155:55]
  wire  _GEN_28197 = next_will_commit_0 & next_will_commit_1 ? _GEN_28004 : _GEN_28132; // @[rob.scala 155:55]
  wire  _GEN_28198 = next_will_commit_0 & next_will_commit_1 ? _GEN_28005 : _GEN_28133; // @[rob.scala 155:55]
  wire  _GEN_28199 = next_will_commit_0 & next_will_commit_1 ? _GEN_28006 : _GEN_28134; // @[rob.scala 155:55]
  wire  _GEN_28200 = next_will_commit_0 & next_will_commit_1 ? _GEN_28007 : _GEN_28135; // @[rob.scala 155:55]
  wire  _GEN_28201 = next_will_commit_0 & next_will_commit_1 ? _GEN_28008 : _GEN_28136; // @[rob.scala 155:55]
  wire  _GEN_28202 = next_will_commit_0 & next_will_commit_1 ? _GEN_28009 : _GEN_28137; // @[rob.scala 155:55]
  wire  _GEN_28203 = next_will_commit_0 & next_will_commit_1 ? _GEN_28010 : _GEN_28138; // @[rob.scala 155:55]
  wire  _GEN_28204 = next_will_commit_0 & next_will_commit_1 ? _GEN_28011 : _GEN_28139; // @[rob.scala 155:55]
  wire  _GEN_28205 = next_will_commit_0 & next_will_commit_1 ? _GEN_28012 : _GEN_28140; // @[rob.scala 155:55]
  wire  _GEN_28206 = next_will_commit_0 & next_will_commit_1 ? _GEN_28013 : _GEN_28141; // @[rob.scala 155:55]
  wire  _GEN_28207 = next_will_commit_0 & next_will_commit_1 ? _GEN_28014 : _GEN_28142; // @[rob.scala 155:55]
  wire  _GEN_28208 = next_will_commit_0 & next_will_commit_1 ? _GEN_28015 : _GEN_28143; // @[rob.scala 155:55]
  wire  _GEN_28209 = next_will_commit_0 & next_will_commit_1 ? _GEN_28016 : _GEN_28144; // @[rob.scala 155:55]
  wire  _GEN_28210 = next_will_commit_0 & next_will_commit_1 ? _GEN_28017 : _GEN_28145; // @[rob.scala 155:55]
  wire  _GEN_28211 = next_will_commit_0 & next_will_commit_1 ? _GEN_28018 : _GEN_28146; // @[rob.scala 155:55]
  wire  _GEN_28212 = next_will_commit_0 & next_will_commit_1 ? _GEN_28019 : _GEN_28147; // @[rob.scala 155:55]
  wire  _GEN_28213 = next_will_commit_0 & next_will_commit_1 ? _GEN_28020 : _GEN_28148; // @[rob.scala 155:55]
  wire  _GEN_28214 = next_will_commit_0 & next_will_commit_1 ? _GEN_28021 : _GEN_28149; // @[rob.scala 155:55]
  wire  _GEN_28215 = next_will_commit_0 & next_will_commit_1 ? _GEN_28022 : _GEN_28150; // @[rob.scala 155:55]
  wire  _GEN_28216 = next_will_commit_0 & next_will_commit_1 ? _GEN_28023 : _GEN_28151; // @[rob.scala 155:55]
  wire  _GEN_28217 = next_will_commit_0 & next_will_commit_1 ? _GEN_28024 : _GEN_28152; // @[rob.scala 155:55]
  wire  _GEN_28218 = next_will_commit_0 & next_will_commit_1 ? _GEN_28025 : _GEN_28153; // @[rob.scala 155:55]
  wire  _GEN_28219 = next_will_commit_0 & next_will_commit_1 ? _GEN_28026 : _GEN_28154; // @[rob.scala 155:55]
  wire  _GEN_28220 = next_will_commit_0 & next_will_commit_1 ? _GEN_28027 : _GEN_28155; // @[rob.scala 155:55]
  wire  _GEN_28221 = next_will_commit_0 & next_will_commit_1 ? _GEN_28028 : _GEN_28156; // @[rob.scala 155:55]
  wire  _GEN_28222 = next_will_commit_0 & next_will_commit_1 ? _GEN_28029 : _GEN_28157; // @[rob.scala 155:55]
  wire  _GEN_28223 = next_will_commit_0 & next_will_commit_1 ? _GEN_28030 : _GEN_28158; // @[rob.scala 155:55]
  wire  _GEN_28224 = next_will_commit_0 & next_will_commit_1 ? _GEN_28031 : _GEN_28159; // @[rob.scala 155:55]
  wire  _GEN_28225 = next_will_commit_0 & next_will_commit_1 ? _GEN_28032 : _GEN_28160; // @[rob.scala 155:55]
  wire  _GEN_28226 = next_will_commit_0 & next_will_commit_1 ? _GEN_28033 : _GEN_28161; // @[rob.scala 155:55]
  wire [6:0] _GEN_28227 = next_will_commit_0 & next_will_commit_1 ? _commit_ptr_T_1 : _GEN_28162; // @[rob.scala 155:55 158:20]
  wire [31:0] _GEN_28292 = _next_will_commit_0_T_5 ? _GEN_25858 : rob_uop_0_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28293 = _next_will_commit_0_T_5 ? _GEN_25859 : rob_uop_1_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28294 = _next_will_commit_0_T_5 ? _GEN_25860 : rob_uop_2_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28295 = _next_will_commit_0_T_5 ? _GEN_25861 : rob_uop_3_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28296 = _next_will_commit_0_T_5 ? _GEN_25862 : rob_uop_4_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28297 = _next_will_commit_0_T_5 ? _GEN_25863 : rob_uop_5_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28298 = _next_will_commit_0_T_5 ? _GEN_25864 : rob_uop_6_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28299 = _next_will_commit_0_T_5 ? _GEN_25865 : rob_uop_7_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28300 = _next_will_commit_0_T_5 ? _GEN_25866 : rob_uop_8_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28301 = _next_will_commit_0_T_5 ? _GEN_25867 : rob_uop_9_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28302 = _next_will_commit_0_T_5 ? _GEN_25868 : rob_uop_10_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28303 = _next_will_commit_0_T_5 ? _GEN_25869 : rob_uop_11_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28304 = _next_will_commit_0_T_5 ? _GEN_25870 : rob_uop_12_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28305 = _next_will_commit_0_T_5 ? _GEN_25871 : rob_uop_13_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28306 = _next_will_commit_0_T_5 ? _GEN_25872 : rob_uop_14_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28307 = _next_will_commit_0_T_5 ? _GEN_25873 : rob_uop_15_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28308 = _next_will_commit_0_T_5 ? _GEN_25874 : rob_uop_16_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28309 = _next_will_commit_0_T_5 ? _GEN_25875 : rob_uop_17_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28310 = _next_will_commit_0_T_5 ? _GEN_25876 : rob_uop_18_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28311 = _next_will_commit_0_T_5 ? _GEN_25877 : rob_uop_19_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28312 = _next_will_commit_0_T_5 ? _GEN_25878 : rob_uop_20_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28313 = _next_will_commit_0_T_5 ? _GEN_25879 : rob_uop_21_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28314 = _next_will_commit_0_T_5 ? _GEN_25880 : rob_uop_22_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28315 = _next_will_commit_0_T_5 ? _GEN_25881 : rob_uop_23_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28316 = _next_will_commit_0_T_5 ? _GEN_25882 : rob_uop_24_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28317 = _next_will_commit_0_T_5 ? _GEN_25883 : rob_uop_25_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28318 = _next_will_commit_0_T_5 ? _GEN_25884 : rob_uop_26_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28319 = _next_will_commit_0_T_5 ? _GEN_25885 : rob_uop_27_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28320 = _next_will_commit_0_T_5 ? _GEN_25886 : rob_uop_28_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28321 = _next_will_commit_0_T_5 ? _GEN_25887 : rob_uop_29_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28322 = _next_will_commit_0_T_5 ? _GEN_25888 : rob_uop_30_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28323 = _next_will_commit_0_T_5 ? _GEN_25889 : rob_uop_31_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28324 = _next_will_commit_0_T_5 ? _GEN_25890 : rob_uop_32_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28325 = _next_will_commit_0_T_5 ? _GEN_25891 : rob_uop_33_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28326 = _next_will_commit_0_T_5 ? _GEN_25892 : rob_uop_34_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28327 = _next_will_commit_0_T_5 ? _GEN_25893 : rob_uop_35_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28328 = _next_will_commit_0_T_5 ? _GEN_25894 : rob_uop_36_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28329 = _next_will_commit_0_T_5 ? _GEN_25895 : rob_uop_37_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28330 = _next_will_commit_0_T_5 ? _GEN_25896 : rob_uop_38_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28331 = _next_will_commit_0_T_5 ? _GEN_25897 : rob_uop_39_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28332 = _next_will_commit_0_T_5 ? _GEN_25898 : rob_uop_40_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28333 = _next_will_commit_0_T_5 ? _GEN_25899 : rob_uop_41_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28334 = _next_will_commit_0_T_5 ? _GEN_25900 : rob_uop_42_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28335 = _next_will_commit_0_T_5 ? _GEN_25901 : rob_uop_43_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28336 = _next_will_commit_0_T_5 ? _GEN_25902 : rob_uop_44_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28337 = _next_will_commit_0_T_5 ? _GEN_25903 : rob_uop_45_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28338 = _next_will_commit_0_T_5 ? _GEN_25904 : rob_uop_46_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28339 = _next_will_commit_0_T_5 ? _GEN_25905 : rob_uop_47_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28340 = _next_will_commit_0_T_5 ? _GEN_25906 : rob_uop_48_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28341 = _next_will_commit_0_T_5 ? _GEN_25907 : rob_uop_49_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28342 = _next_will_commit_0_T_5 ? _GEN_25908 : rob_uop_50_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28343 = _next_will_commit_0_T_5 ? _GEN_25909 : rob_uop_51_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28344 = _next_will_commit_0_T_5 ? _GEN_25910 : rob_uop_52_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28345 = _next_will_commit_0_T_5 ? _GEN_25911 : rob_uop_53_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28346 = _next_will_commit_0_T_5 ? _GEN_25912 : rob_uop_54_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28347 = _next_will_commit_0_T_5 ? _GEN_25913 : rob_uop_55_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28348 = _next_will_commit_0_T_5 ? _GEN_25914 : rob_uop_56_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28349 = _next_will_commit_0_T_5 ? _GEN_25915 : rob_uop_57_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28350 = _next_will_commit_0_T_5 ? _GEN_25916 : rob_uop_58_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28351 = _next_will_commit_0_T_5 ? _GEN_25917 : rob_uop_59_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28352 = _next_will_commit_0_T_5 ? _GEN_25918 : rob_uop_60_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28353 = _next_will_commit_0_T_5 ? _GEN_25919 : rob_uop_61_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28354 = _next_will_commit_0_T_5 ? _GEN_25920 : rob_uop_62_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28355 = _next_will_commit_0_T_5 ? _GEN_25921 : rob_uop_63_pc; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28356 = _next_will_commit_0_T_5 ? _GEN_25922 : rob_uop_0_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28357 = _next_will_commit_0_T_5 ? _GEN_25923 : rob_uop_1_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28358 = _next_will_commit_0_T_5 ? _GEN_25924 : rob_uop_2_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28359 = _next_will_commit_0_T_5 ? _GEN_25925 : rob_uop_3_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28360 = _next_will_commit_0_T_5 ? _GEN_25926 : rob_uop_4_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28361 = _next_will_commit_0_T_5 ? _GEN_25927 : rob_uop_5_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28362 = _next_will_commit_0_T_5 ? _GEN_25928 : rob_uop_6_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28363 = _next_will_commit_0_T_5 ? _GEN_25929 : rob_uop_7_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28364 = _next_will_commit_0_T_5 ? _GEN_25930 : rob_uop_8_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28365 = _next_will_commit_0_T_5 ? _GEN_25931 : rob_uop_9_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28366 = _next_will_commit_0_T_5 ? _GEN_25932 : rob_uop_10_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28367 = _next_will_commit_0_T_5 ? _GEN_25933 : rob_uop_11_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28368 = _next_will_commit_0_T_5 ? _GEN_25934 : rob_uop_12_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28369 = _next_will_commit_0_T_5 ? _GEN_25935 : rob_uop_13_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28370 = _next_will_commit_0_T_5 ? _GEN_25936 : rob_uop_14_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28371 = _next_will_commit_0_T_5 ? _GEN_25937 : rob_uop_15_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28372 = _next_will_commit_0_T_5 ? _GEN_25938 : rob_uop_16_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28373 = _next_will_commit_0_T_5 ? _GEN_25939 : rob_uop_17_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28374 = _next_will_commit_0_T_5 ? _GEN_25940 : rob_uop_18_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28375 = _next_will_commit_0_T_5 ? _GEN_25941 : rob_uop_19_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28376 = _next_will_commit_0_T_5 ? _GEN_25942 : rob_uop_20_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28377 = _next_will_commit_0_T_5 ? _GEN_25943 : rob_uop_21_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28378 = _next_will_commit_0_T_5 ? _GEN_25944 : rob_uop_22_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28379 = _next_will_commit_0_T_5 ? _GEN_25945 : rob_uop_23_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28380 = _next_will_commit_0_T_5 ? _GEN_25946 : rob_uop_24_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28381 = _next_will_commit_0_T_5 ? _GEN_25947 : rob_uop_25_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28382 = _next_will_commit_0_T_5 ? _GEN_25948 : rob_uop_26_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28383 = _next_will_commit_0_T_5 ? _GEN_25949 : rob_uop_27_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28384 = _next_will_commit_0_T_5 ? _GEN_25950 : rob_uop_28_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28385 = _next_will_commit_0_T_5 ? _GEN_25951 : rob_uop_29_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28386 = _next_will_commit_0_T_5 ? _GEN_25952 : rob_uop_30_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28387 = _next_will_commit_0_T_5 ? _GEN_25953 : rob_uop_31_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28388 = _next_will_commit_0_T_5 ? _GEN_25954 : rob_uop_32_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28389 = _next_will_commit_0_T_5 ? _GEN_25955 : rob_uop_33_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28390 = _next_will_commit_0_T_5 ? _GEN_25956 : rob_uop_34_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28391 = _next_will_commit_0_T_5 ? _GEN_25957 : rob_uop_35_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28392 = _next_will_commit_0_T_5 ? _GEN_25958 : rob_uop_36_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28393 = _next_will_commit_0_T_5 ? _GEN_25959 : rob_uop_37_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28394 = _next_will_commit_0_T_5 ? _GEN_25960 : rob_uop_38_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28395 = _next_will_commit_0_T_5 ? _GEN_25961 : rob_uop_39_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28396 = _next_will_commit_0_T_5 ? _GEN_25962 : rob_uop_40_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28397 = _next_will_commit_0_T_5 ? _GEN_25963 : rob_uop_41_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28398 = _next_will_commit_0_T_5 ? _GEN_25964 : rob_uop_42_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28399 = _next_will_commit_0_T_5 ? _GEN_25965 : rob_uop_43_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28400 = _next_will_commit_0_T_5 ? _GEN_25966 : rob_uop_44_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28401 = _next_will_commit_0_T_5 ? _GEN_25967 : rob_uop_45_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28402 = _next_will_commit_0_T_5 ? _GEN_25968 : rob_uop_46_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28403 = _next_will_commit_0_T_5 ? _GEN_25969 : rob_uop_47_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28404 = _next_will_commit_0_T_5 ? _GEN_25970 : rob_uop_48_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28405 = _next_will_commit_0_T_5 ? _GEN_25971 : rob_uop_49_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28406 = _next_will_commit_0_T_5 ? _GEN_25972 : rob_uop_50_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28407 = _next_will_commit_0_T_5 ? _GEN_25973 : rob_uop_51_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28408 = _next_will_commit_0_T_5 ? _GEN_25974 : rob_uop_52_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28409 = _next_will_commit_0_T_5 ? _GEN_25975 : rob_uop_53_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28410 = _next_will_commit_0_T_5 ? _GEN_25976 : rob_uop_54_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28411 = _next_will_commit_0_T_5 ? _GEN_25977 : rob_uop_55_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28412 = _next_will_commit_0_T_5 ? _GEN_25978 : rob_uop_56_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28413 = _next_will_commit_0_T_5 ? _GEN_25979 : rob_uop_57_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28414 = _next_will_commit_0_T_5 ? _GEN_25980 : rob_uop_58_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28415 = _next_will_commit_0_T_5 ? _GEN_25981 : rob_uop_59_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28416 = _next_will_commit_0_T_5 ? _GEN_25982 : rob_uop_60_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28417 = _next_will_commit_0_T_5 ? _GEN_25983 : rob_uop_61_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28418 = _next_will_commit_0_T_5 ? _GEN_25984 : rob_uop_62_inst; // @[rob.scala 123:38 82:26]
  wire [31:0] _GEN_28419 = _next_will_commit_0_T_5 ? _GEN_25985 : rob_uop_63_inst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28420 = _next_will_commit_0_T_5 ? _GEN_25986 : rob_uop_0_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28421 = _next_will_commit_0_T_5 ? _GEN_25987 : rob_uop_1_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28422 = _next_will_commit_0_T_5 ? _GEN_25988 : rob_uop_2_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28423 = _next_will_commit_0_T_5 ? _GEN_25989 : rob_uop_3_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28424 = _next_will_commit_0_T_5 ? _GEN_25990 : rob_uop_4_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28425 = _next_will_commit_0_T_5 ? _GEN_25991 : rob_uop_5_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28426 = _next_will_commit_0_T_5 ? _GEN_25992 : rob_uop_6_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28427 = _next_will_commit_0_T_5 ? _GEN_25993 : rob_uop_7_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28428 = _next_will_commit_0_T_5 ? _GEN_25994 : rob_uop_8_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28429 = _next_will_commit_0_T_5 ? _GEN_25995 : rob_uop_9_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28430 = _next_will_commit_0_T_5 ? _GEN_25996 : rob_uop_10_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28431 = _next_will_commit_0_T_5 ? _GEN_25997 : rob_uop_11_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28432 = _next_will_commit_0_T_5 ? _GEN_25998 : rob_uop_12_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28433 = _next_will_commit_0_T_5 ? _GEN_25999 : rob_uop_13_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28434 = _next_will_commit_0_T_5 ? _GEN_26000 : rob_uop_14_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28435 = _next_will_commit_0_T_5 ? _GEN_26001 : rob_uop_15_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28436 = _next_will_commit_0_T_5 ? _GEN_26002 : rob_uop_16_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28437 = _next_will_commit_0_T_5 ? _GEN_26003 : rob_uop_17_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28438 = _next_will_commit_0_T_5 ? _GEN_26004 : rob_uop_18_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28439 = _next_will_commit_0_T_5 ? _GEN_26005 : rob_uop_19_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28440 = _next_will_commit_0_T_5 ? _GEN_26006 : rob_uop_20_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28441 = _next_will_commit_0_T_5 ? _GEN_26007 : rob_uop_21_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28442 = _next_will_commit_0_T_5 ? _GEN_26008 : rob_uop_22_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28443 = _next_will_commit_0_T_5 ? _GEN_26009 : rob_uop_23_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28444 = _next_will_commit_0_T_5 ? _GEN_26010 : rob_uop_24_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28445 = _next_will_commit_0_T_5 ? _GEN_26011 : rob_uop_25_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28446 = _next_will_commit_0_T_5 ? _GEN_26012 : rob_uop_26_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28447 = _next_will_commit_0_T_5 ? _GEN_26013 : rob_uop_27_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28448 = _next_will_commit_0_T_5 ? _GEN_26014 : rob_uop_28_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28449 = _next_will_commit_0_T_5 ? _GEN_26015 : rob_uop_29_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28450 = _next_will_commit_0_T_5 ? _GEN_26016 : rob_uop_30_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28451 = _next_will_commit_0_T_5 ? _GEN_26017 : rob_uop_31_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28452 = _next_will_commit_0_T_5 ? _GEN_26018 : rob_uop_32_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28453 = _next_will_commit_0_T_5 ? _GEN_26019 : rob_uop_33_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28454 = _next_will_commit_0_T_5 ? _GEN_26020 : rob_uop_34_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28455 = _next_will_commit_0_T_5 ? _GEN_26021 : rob_uop_35_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28456 = _next_will_commit_0_T_5 ? _GEN_26022 : rob_uop_36_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28457 = _next_will_commit_0_T_5 ? _GEN_26023 : rob_uop_37_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28458 = _next_will_commit_0_T_5 ? _GEN_26024 : rob_uop_38_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28459 = _next_will_commit_0_T_5 ? _GEN_26025 : rob_uop_39_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28460 = _next_will_commit_0_T_5 ? _GEN_26026 : rob_uop_40_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28461 = _next_will_commit_0_T_5 ? _GEN_26027 : rob_uop_41_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28462 = _next_will_commit_0_T_5 ? _GEN_26028 : rob_uop_42_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28463 = _next_will_commit_0_T_5 ? _GEN_26029 : rob_uop_43_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28464 = _next_will_commit_0_T_5 ? _GEN_26030 : rob_uop_44_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28465 = _next_will_commit_0_T_5 ? _GEN_26031 : rob_uop_45_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28466 = _next_will_commit_0_T_5 ? _GEN_26032 : rob_uop_46_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28467 = _next_will_commit_0_T_5 ? _GEN_26033 : rob_uop_47_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28468 = _next_will_commit_0_T_5 ? _GEN_26034 : rob_uop_48_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28469 = _next_will_commit_0_T_5 ? _GEN_26035 : rob_uop_49_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28470 = _next_will_commit_0_T_5 ? _GEN_26036 : rob_uop_50_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28471 = _next_will_commit_0_T_5 ? _GEN_26037 : rob_uop_51_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28472 = _next_will_commit_0_T_5 ? _GEN_26038 : rob_uop_52_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28473 = _next_will_commit_0_T_5 ? _GEN_26039 : rob_uop_53_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28474 = _next_will_commit_0_T_5 ? _GEN_26040 : rob_uop_54_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28475 = _next_will_commit_0_T_5 ? _GEN_26041 : rob_uop_55_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28476 = _next_will_commit_0_T_5 ? _GEN_26042 : rob_uop_56_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28477 = _next_will_commit_0_T_5 ? _GEN_26043 : rob_uop_57_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28478 = _next_will_commit_0_T_5 ? _GEN_26044 : rob_uop_58_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28479 = _next_will_commit_0_T_5 ? _GEN_26045 : rob_uop_59_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28480 = _next_will_commit_0_T_5 ? _GEN_26046 : rob_uop_60_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28481 = _next_will_commit_0_T_5 ? _GEN_26047 : rob_uop_61_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28482 = _next_will_commit_0_T_5 ? _GEN_26048 : rob_uop_62_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28483 = _next_will_commit_0_T_5 ? _GEN_26049 : rob_uop_63_func_code; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28804 = _next_will_commit_0_T_5 ? _GEN_26370 : rob_uop_0_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28805 = _next_will_commit_0_T_5 ? _GEN_26371 : rob_uop_1_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28806 = _next_will_commit_0_T_5 ? _GEN_26372 : rob_uop_2_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28807 = _next_will_commit_0_T_5 ? _GEN_26373 : rob_uop_3_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28808 = _next_will_commit_0_T_5 ? _GEN_26374 : rob_uop_4_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28809 = _next_will_commit_0_T_5 ? _GEN_26375 : rob_uop_5_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28810 = _next_will_commit_0_T_5 ? _GEN_26376 : rob_uop_6_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28811 = _next_will_commit_0_T_5 ? _GEN_26377 : rob_uop_7_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28812 = _next_will_commit_0_T_5 ? _GEN_26378 : rob_uop_8_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28813 = _next_will_commit_0_T_5 ? _GEN_26379 : rob_uop_9_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28814 = _next_will_commit_0_T_5 ? _GEN_26380 : rob_uop_10_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28815 = _next_will_commit_0_T_5 ? _GEN_26381 : rob_uop_11_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28816 = _next_will_commit_0_T_5 ? _GEN_26382 : rob_uop_12_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28817 = _next_will_commit_0_T_5 ? _GEN_26383 : rob_uop_13_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28818 = _next_will_commit_0_T_5 ? _GEN_26384 : rob_uop_14_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28819 = _next_will_commit_0_T_5 ? _GEN_26385 : rob_uop_15_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28820 = _next_will_commit_0_T_5 ? _GEN_26386 : rob_uop_16_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28821 = _next_will_commit_0_T_5 ? _GEN_26387 : rob_uop_17_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28822 = _next_will_commit_0_T_5 ? _GEN_26388 : rob_uop_18_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28823 = _next_will_commit_0_T_5 ? _GEN_26389 : rob_uop_19_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28824 = _next_will_commit_0_T_5 ? _GEN_26390 : rob_uop_20_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28825 = _next_will_commit_0_T_5 ? _GEN_26391 : rob_uop_21_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28826 = _next_will_commit_0_T_5 ? _GEN_26392 : rob_uop_22_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28827 = _next_will_commit_0_T_5 ? _GEN_26393 : rob_uop_23_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28828 = _next_will_commit_0_T_5 ? _GEN_26394 : rob_uop_24_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28829 = _next_will_commit_0_T_5 ? _GEN_26395 : rob_uop_25_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28830 = _next_will_commit_0_T_5 ? _GEN_26396 : rob_uop_26_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28831 = _next_will_commit_0_T_5 ? _GEN_26397 : rob_uop_27_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28832 = _next_will_commit_0_T_5 ? _GEN_26398 : rob_uop_28_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28833 = _next_will_commit_0_T_5 ? _GEN_26399 : rob_uop_29_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28834 = _next_will_commit_0_T_5 ? _GEN_26400 : rob_uop_30_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28835 = _next_will_commit_0_T_5 ? _GEN_26401 : rob_uop_31_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28836 = _next_will_commit_0_T_5 ? _GEN_26402 : rob_uop_32_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28837 = _next_will_commit_0_T_5 ? _GEN_26403 : rob_uop_33_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28838 = _next_will_commit_0_T_5 ? _GEN_26404 : rob_uop_34_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28839 = _next_will_commit_0_T_5 ? _GEN_26405 : rob_uop_35_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28840 = _next_will_commit_0_T_5 ? _GEN_26406 : rob_uop_36_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28841 = _next_will_commit_0_T_5 ? _GEN_26407 : rob_uop_37_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28842 = _next_will_commit_0_T_5 ? _GEN_26408 : rob_uop_38_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28843 = _next_will_commit_0_T_5 ? _GEN_26409 : rob_uop_39_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28844 = _next_will_commit_0_T_5 ? _GEN_26410 : rob_uop_40_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28845 = _next_will_commit_0_T_5 ? _GEN_26411 : rob_uop_41_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28846 = _next_will_commit_0_T_5 ? _GEN_26412 : rob_uop_42_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28847 = _next_will_commit_0_T_5 ? _GEN_26413 : rob_uop_43_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28848 = _next_will_commit_0_T_5 ? _GEN_26414 : rob_uop_44_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28849 = _next_will_commit_0_T_5 ? _GEN_26415 : rob_uop_45_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28850 = _next_will_commit_0_T_5 ? _GEN_26416 : rob_uop_46_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28851 = _next_will_commit_0_T_5 ? _GEN_26417 : rob_uop_47_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28852 = _next_will_commit_0_T_5 ? _GEN_26418 : rob_uop_48_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28853 = _next_will_commit_0_T_5 ? _GEN_26419 : rob_uop_49_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28854 = _next_will_commit_0_T_5 ? _GEN_26420 : rob_uop_50_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28855 = _next_will_commit_0_T_5 ? _GEN_26421 : rob_uop_51_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28856 = _next_will_commit_0_T_5 ? _GEN_26422 : rob_uop_52_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28857 = _next_will_commit_0_T_5 ? _GEN_26423 : rob_uop_53_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28858 = _next_will_commit_0_T_5 ? _GEN_26424 : rob_uop_54_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28859 = _next_will_commit_0_T_5 ? _GEN_26425 : rob_uop_55_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28860 = _next_will_commit_0_T_5 ? _GEN_26426 : rob_uop_56_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28861 = _next_will_commit_0_T_5 ? _GEN_26427 : rob_uop_57_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28862 = _next_will_commit_0_T_5 ? _GEN_26428 : rob_uop_58_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28863 = _next_will_commit_0_T_5 ? _GEN_26429 : rob_uop_59_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28864 = _next_will_commit_0_T_5 ? _GEN_26430 : rob_uop_60_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28865 = _next_will_commit_0_T_5 ? _GEN_26431 : rob_uop_61_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28866 = _next_will_commit_0_T_5 ? _GEN_26432 : rob_uop_62_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28867 = _next_will_commit_0_T_5 ? _GEN_26433 : rob_uop_63_phy_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28868 = _next_will_commit_0_T_5 ? _GEN_26434 : rob_uop_0_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28869 = _next_will_commit_0_T_5 ? _GEN_26435 : rob_uop_1_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28870 = _next_will_commit_0_T_5 ? _GEN_26436 : rob_uop_2_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28871 = _next_will_commit_0_T_5 ? _GEN_26437 : rob_uop_3_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28872 = _next_will_commit_0_T_5 ? _GEN_26438 : rob_uop_4_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28873 = _next_will_commit_0_T_5 ? _GEN_26439 : rob_uop_5_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28874 = _next_will_commit_0_T_5 ? _GEN_26440 : rob_uop_6_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28875 = _next_will_commit_0_T_5 ? _GEN_26441 : rob_uop_7_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28876 = _next_will_commit_0_T_5 ? _GEN_26442 : rob_uop_8_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28877 = _next_will_commit_0_T_5 ? _GEN_26443 : rob_uop_9_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28878 = _next_will_commit_0_T_5 ? _GEN_26444 : rob_uop_10_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28879 = _next_will_commit_0_T_5 ? _GEN_26445 : rob_uop_11_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28880 = _next_will_commit_0_T_5 ? _GEN_26446 : rob_uop_12_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28881 = _next_will_commit_0_T_5 ? _GEN_26447 : rob_uop_13_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28882 = _next_will_commit_0_T_5 ? _GEN_26448 : rob_uop_14_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28883 = _next_will_commit_0_T_5 ? _GEN_26449 : rob_uop_15_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28884 = _next_will_commit_0_T_5 ? _GEN_26450 : rob_uop_16_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28885 = _next_will_commit_0_T_5 ? _GEN_26451 : rob_uop_17_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28886 = _next_will_commit_0_T_5 ? _GEN_26452 : rob_uop_18_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28887 = _next_will_commit_0_T_5 ? _GEN_26453 : rob_uop_19_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28888 = _next_will_commit_0_T_5 ? _GEN_26454 : rob_uop_20_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28889 = _next_will_commit_0_T_5 ? _GEN_26455 : rob_uop_21_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28890 = _next_will_commit_0_T_5 ? _GEN_26456 : rob_uop_22_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28891 = _next_will_commit_0_T_5 ? _GEN_26457 : rob_uop_23_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28892 = _next_will_commit_0_T_5 ? _GEN_26458 : rob_uop_24_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28893 = _next_will_commit_0_T_5 ? _GEN_26459 : rob_uop_25_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28894 = _next_will_commit_0_T_5 ? _GEN_26460 : rob_uop_26_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28895 = _next_will_commit_0_T_5 ? _GEN_26461 : rob_uop_27_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28896 = _next_will_commit_0_T_5 ? _GEN_26462 : rob_uop_28_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28897 = _next_will_commit_0_T_5 ? _GEN_26463 : rob_uop_29_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28898 = _next_will_commit_0_T_5 ? _GEN_26464 : rob_uop_30_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28899 = _next_will_commit_0_T_5 ? _GEN_26465 : rob_uop_31_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28900 = _next_will_commit_0_T_5 ? _GEN_26466 : rob_uop_32_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28901 = _next_will_commit_0_T_5 ? _GEN_26467 : rob_uop_33_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28902 = _next_will_commit_0_T_5 ? _GEN_26468 : rob_uop_34_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28903 = _next_will_commit_0_T_5 ? _GEN_26469 : rob_uop_35_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28904 = _next_will_commit_0_T_5 ? _GEN_26470 : rob_uop_36_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28905 = _next_will_commit_0_T_5 ? _GEN_26471 : rob_uop_37_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28906 = _next_will_commit_0_T_5 ? _GEN_26472 : rob_uop_38_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28907 = _next_will_commit_0_T_5 ? _GEN_26473 : rob_uop_39_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28908 = _next_will_commit_0_T_5 ? _GEN_26474 : rob_uop_40_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28909 = _next_will_commit_0_T_5 ? _GEN_26475 : rob_uop_41_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28910 = _next_will_commit_0_T_5 ? _GEN_26476 : rob_uop_42_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28911 = _next_will_commit_0_T_5 ? _GEN_26477 : rob_uop_43_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28912 = _next_will_commit_0_T_5 ? _GEN_26478 : rob_uop_44_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28913 = _next_will_commit_0_T_5 ? _GEN_26479 : rob_uop_45_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28914 = _next_will_commit_0_T_5 ? _GEN_26480 : rob_uop_46_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28915 = _next_will_commit_0_T_5 ? _GEN_26481 : rob_uop_47_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28916 = _next_will_commit_0_T_5 ? _GEN_26482 : rob_uop_48_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28917 = _next_will_commit_0_T_5 ? _GEN_26483 : rob_uop_49_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28918 = _next_will_commit_0_T_5 ? _GEN_26484 : rob_uop_50_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28919 = _next_will_commit_0_T_5 ? _GEN_26485 : rob_uop_51_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28920 = _next_will_commit_0_T_5 ? _GEN_26486 : rob_uop_52_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28921 = _next_will_commit_0_T_5 ? _GEN_26487 : rob_uop_53_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28922 = _next_will_commit_0_T_5 ? _GEN_26488 : rob_uop_54_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28923 = _next_will_commit_0_T_5 ? _GEN_26489 : rob_uop_55_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28924 = _next_will_commit_0_T_5 ? _GEN_26490 : rob_uop_56_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28925 = _next_will_commit_0_T_5 ? _GEN_26491 : rob_uop_57_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28926 = _next_will_commit_0_T_5 ? _GEN_26492 : rob_uop_58_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28927 = _next_will_commit_0_T_5 ? _GEN_26493 : rob_uop_59_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28928 = _next_will_commit_0_T_5 ? _GEN_26494 : rob_uop_60_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28929 = _next_will_commit_0_T_5 ? _GEN_26495 : rob_uop_61_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28930 = _next_will_commit_0_T_5 ? _GEN_26496 : rob_uop_62_stale_dst; // @[rob.scala 123:38 82:26]
  wire [6:0] _GEN_28931 = _next_will_commit_0_T_5 ? _GEN_26497 : rob_uop_63_stale_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28932 = _next_will_commit_0_T_5 ? _GEN_26498 : rob_uop_0_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28933 = _next_will_commit_0_T_5 ? _GEN_26499 : rob_uop_1_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28934 = _next_will_commit_0_T_5 ? _GEN_26500 : rob_uop_2_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28935 = _next_will_commit_0_T_5 ? _GEN_26501 : rob_uop_3_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28936 = _next_will_commit_0_T_5 ? _GEN_26502 : rob_uop_4_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28937 = _next_will_commit_0_T_5 ? _GEN_26503 : rob_uop_5_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28938 = _next_will_commit_0_T_5 ? _GEN_26504 : rob_uop_6_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28939 = _next_will_commit_0_T_5 ? _GEN_26505 : rob_uop_7_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28940 = _next_will_commit_0_T_5 ? _GEN_26506 : rob_uop_8_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28941 = _next_will_commit_0_T_5 ? _GEN_26507 : rob_uop_9_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28942 = _next_will_commit_0_T_5 ? _GEN_26508 : rob_uop_10_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28943 = _next_will_commit_0_T_5 ? _GEN_26509 : rob_uop_11_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28944 = _next_will_commit_0_T_5 ? _GEN_26510 : rob_uop_12_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28945 = _next_will_commit_0_T_5 ? _GEN_26511 : rob_uop_13_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28946 = _next_will_commit_0_T_5 ? _GEN_26512 : rob_uop_14_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28947 = _next_will_commit_0_T_5 ? _GEN_26513 : rob_uop_15_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28948 = _next_will_commit_0_T_5 ? _GEN_26514 : rob_uop_16_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28949 = _next_will_commit_0_T_5 ? _GEN_26515 : rob_uop_17_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28950 = _next_will_commit_0_T_5 ? _GEN_26516 : rob_uop_18_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28951 = _next_will_commit_0_T_5 ? _GEN_26517 : rob_uop_19_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28952 = _next_will_commit_0_T_5 ? _GEN_26518 : rob_uop_20_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28953 = _next_will_commit_0_T_5 ? _GEN_26519 : rob_uop_21_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28954 = _next_will_commit_0_T_5 ? _GEN_26520 : rob_uop_22_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28955 = _next_will_commit_0_T_5 ? _GEN_26521 : rob_uop_23_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28956 = _next_will_commit_0_T_5 ? _GEN_26522 : rob_uop_24_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28957 = _next_will_commit_0_T_5 ? _GEN_26523 : rob_uop_25_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28958 = _next_will_commit_0_T_5 ? _GEN_26524 : rob_uop_26_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28959 = _next_will_commit_0_T_5 ? _GEN_26525 : rob_uop_27_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28960 = _next_will_commit_0_T_5 ? _GEN_26526 : rob_uop_28_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28961 = _next_will_commit_0_T_5 ? _GEN_26527 : rob_uop_29_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28962 = _next_will_commit_0_T_5 ? _GEN_26528 : rob_uop_30_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28963 = _next_will_commit_0_T_5 ? _GEN_26529 : rob_uop_31_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28964 = _next_will_commit_0_T_5 ? _GEN_26530 : rob_uop_32_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28965 = _next_will_commit_0_T_5 ? _GEN_26531 : rob_uop_33_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28966 = _next_will_commit_0_T_5 ? _GEN_26532 : rob_uop_34_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28967 = _next_will_commit_0_T_5 ? _GEN_26533 : rob_uop_35_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28968 = _next_will_commit_0_T_5 ? _GEN_26534 : rob_uop_36_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28969 = _next_will_commit_0_T_5 ? _GEN_26535 : rob_uop_37_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28970 = _next_will_commit_0_T_5 ? _GEN_26536 : rob_uop_38_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28971 = _next_will_commit_0_T_5 ? _GEN_26537 : rob_uop_39_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28972 = _next_will_commit_0_T_5 ? _GEN_26538 : rob_uop_40_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28973 = _next_will_commit_0_T_5 ? _GEN_26539 : rob_uop_41_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28974 = _next_will_commit_0_T_5 ? _GEN_26540 : rob_uop_42_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28975 = _next_will_commit_0_T_5 ? _GEN_26541 : rob_uop_43_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28976 = _next_will_commit_0_T_5 ? _GEN_26542 : rob_uop_44_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28977 = _next_will_commit_0_T_5 ? _GEN_26543 : rob_uop_45_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28978 = _next_will_commit_0_T_5 ? _GEN_26544 : rob_uop_46_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28979 = _next_will_commit_0_T_5 ? _GEN_26545 : rob_uop_47_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28980 = _next_will_commit_0_T_5 ? _GEN_26546 : rob_uop_48_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28981 = _next_will_commit_0_T_5 ? _GEN_26547 : rob_uop_49_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28982 = _next_will_commit_0_T_5 ? _GEN_26548 : rob_uop_50_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28983 = _next_will_commit_0_T_5 ? _GEN_26549 : rob_uop_51_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28984 = _next_will_commit_0_T_5 ? _GEN_26550 : rob_uop_52_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28985 = _next_will_commit_0_T_5 ? _GEN_26551 : rob_uop_53_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28986 = _next_will_commit_0_T_5 ? _GEN_26552 : rob_uop_54_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28987 = _next_will_commit_0_T_5 ? _GEN_26553 : rob_uop_55_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28988 = _next_will_commit_0_T_5 ? _GEN_26554 : rob_uop_56_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28989 = _next_will_commit_0_T_5 ? _GEN_26555 : rob_uop_57_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28990 = _next_will_commit_0_T_5 ? _GEN_26556 : rob_uop_58_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28991 = _next_will_commit_0_T_5 ? _GEN_26557 : rob_uop_59_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28992 = _next_will_commit_0_T_5 ? _GEN_26558 : rob_uop_60_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28993 = _next_will_commit_0_T_5 ? _GEN_26559 : rob_uop_61_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28994 = _next_will_commit_0_T_5 ? _GEN_26560 : rob_uop_62_arch_dst; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_28995 = _next_will_commit_0_T_5 ? _GEN_26561 : rob_uop_63_arch_dst; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29636 = _next_will_commit_0_T_5 ? _GEN_27202 : rob_uop_0_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29637 = _next_will_commit_0_T_5 ? _GEN_27203 : rob_uop_1_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29638 = _next_will_commit_0_T_5 ? _GEN_27204 : rob_uop_2_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29639 = _next_will_commit_0_T_5 ? _GEN_27205 : rob_uop_3_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29640 = _next_will_commit_0_T_5 ? _GEN_27206 : rob_uop_4_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29641 = _next_will_commit_0_T_5 ? _GEN_27207 : rob_uop_5_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29642 = _next_will_commit_0_T_5 ? _GEN_27208 : rob_uop_6_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29643 = _next_will_commit_0_T_5 ? _GEN_27209 : rob_uop_7_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29644 = _next_will_commit_0_T_5 ? _GEN_27210 : rob_uop_8_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29645 = _next_will_commit_0_T_5 ? _GEN_27211 : rob_uop_9_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29646 = _next_will_commit_0_T_5 ? _GEN_27212 : rob_uop_10_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29647 = _next_will_commit_0_T_5 ? _GEN_27213 : rob_uop_11_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29648 = _next_will_commit_0_T_5 ? _GEN_27214 : rob_uop_12_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29649 = _next_will_commit_0_T_5 ? _GEN_27215 : rob_uop_13_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29650 = _next_will_commit_0_T_5 ? _GEN_27216 : rob_uop_14_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29651 = _next_will_commit_0_T_5 ? _GEN_27217 : rob_uop_15_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29652 = _next_will_commit_0_T_5 ? _GEN_27218 : rob_uop_16_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29653 = _next_will_commit_0_T_5 ? _GEN_27219 : rob_uop_17_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29654 = _next_will_commit_0_T_5 ? _GEN_27220 : rob_uop_18_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29655 = _next_will_commit_0_T_5 ? _GEN_27221 : rob_uop_19_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29656 = _next_will_commit_0_T_5 ? _GEN_27222 : rob_uop_20_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29657 = _next_will_commit_0_T_5 ? _GEN_27223 : rob_uop_21_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29658 = _next_will_commit_0_T_5 ? _GEN_27224 : rob_uop_22_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29659 = _next_will_commit_0_T_5 ? _GEN_27225 : rob_uop_23_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29660 = _next_will_commit_0_T_5 ? _GEN_27226 : rob_uop_24_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29661 = _next_will_commit_0_T_5 ? _GEN_27227 : rob_uop_25_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29662 = _next_will_commit_0_T_5 ? _GEN_27228 : rob_uop_26_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29663 = _next_will_commit_0_T_5 ? _GEN_27229 : rob_uop_27_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29664 = _next_will_commit_0_T_5 ? _GEN_27230 : rob_uop_28_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29665 = _next_will_commit_0_T_5 ? _GEN_27231 : rob_uop_29_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29666 = _next_will_commit_0_T_5 ? _GEN_27232 : rob_uop_30_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29667 = _next_will_commit_0_T_5 ? _GEN_27233 : rob_uop_31_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29668 = _next_will_commit_0_T_5 ? _GEN_27234 : rob_uop_32_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29669 = _next_will_commit_0_T_5 ? _GEN_27235 : rob_uop_33_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29670 = _next_will_commit_0_T_5 ? _GEN_27236 : rob_uop_34_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29671 = _next_will_commit_0_T_5 ? _GEN_27237 : rob_uop_35_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29672 = _next_will_commit_0_T_5 ? _GEN_27238 : rob_uop_36_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29673 = _next_will_commit_0_T_5 ? _GEN_27239 : rob_uop_37_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29674 = _next_will_commit_0_T_5 ? _GEN_27240 : rob_uop_38_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29675 = _next_will_commit_0_T_5 ? _GEN_27241 : rob_uop_39_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29676 = _next_will_commit_0_T_5 ? _GEN_27242 : rob_uop_40_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29677 = _next_will_commit_0_T_5 ? _GEN_27243 : rob_uop_41_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29678 = _next_will_commit_0_T_5 ? _GEN_27244 : rob_uop_42_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29679 = _next_will_commit_0_T_5 ? _GEN_27245 : rob_uop_43_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29680 = _next_will_commit_0_T_5 ? _GEN_27246 : rob_uop_44_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29681 = _next_will_commit_0_T_5 ? _GEN_27247 : rob_uop_45_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29682 = _next_will_commit_0_T_5 ? _GEN_27248 : rob_uop_46_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29683 = _next_will_commit_0_T_5 ? _GEN_27249 : rob_uop_47_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29684 = _next_will_commit_0_T_5 ? _GEN_27250 : rob_uop_48_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29685 = _next_will_commit_0_T_5 ? _GEN_27251 : rob_uop_49_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29686 = _next_will_commit_0_T_5 ? _GEN_27252 : rob_uop_50_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29687 = _next_will_commit_0_T_5 ? _GEN_27253 : rob_uop_51_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29688 = _next_will_commit_0_T_5 ? _GEN_27254 : rob_uop_52_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29689 = _next_will_commit_0_T_5 ? _GEN_27255 : rob_uop_53_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29690 = _next_will_commit_0_T_5 ? _GEN_27256 : rob_uop_54_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29691 = _next_will_commit_0_T_5 ? _GEN_27257 : rob_uop_55_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29692 = _next_will_commit_0_T_5 ? _GEN_27258 : rob_uop_56_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29693 = _next_will_commit_0_T_5 ? _GEN_27259 : rob_uop_57_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29694 = _next_will_commit_0_T_5 ? _GEN_27260 : rob_uop_58_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29695 = _next_will_commit_0_T_5 ? _GEN_27261 : rob_uop_59_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29696 = _next_will_commit_0_T_5 ? _GEN_27262 : rob_uop_60_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29697 = _next_will_commit_0_T_5 ? _GEN_27263 : rob_uop_61_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29698 = _next_will_commit_0_T_5 ? _GEN_27264 : rob_uop_62_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29699 = _next_will_commit_0_T_5 ? _GEN_27265 : rob_uop_63_dst_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29700 = _next_will_commit_0_T_5 ? _GEN_27266 : rob_uop_0_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29701 = _next_will_commit_0_T_5 ? _GEN_27267 : rob_uop_1_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29702 = _next_will_commit_0_T_5 ? _GEN_27268 : rob_uop_2_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29703 = _next_will_commit_0_T_5 ? _GEN_27269 : rob_uop_3_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29704 = _next_will_commit_0_T_5 ? _GEN_27270 : rob_uop_4_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29705 = _next_will_commit_0_T_5 ? _GEN_27271 : rob_uop_5_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29706 = _next_will_commit_0_T_5 ? _GEN_27272 : rob_uop_6_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29707 = _next_will_commit_0_T_5 ? _GEN_27273 : rob_uop_7_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29708 = _next_will_commit_0_T_5 ? _GEN_27274 : rob_uop_8_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29709 = _next_will_commit_0_T_5 ? _GEN_27275 : rob_uop_9_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29710 = _next_will_commit_0_T_5 ? _GEN_27276 : rob_uop_10_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29711 = _next_will_commit_0_T_5 ? _GEN_27277 : rob_uop_11_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29712 = _next_will_commit_0_T_5 ? _GEN_27278 : rob_uop_12_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29713 = _next_will_commit_0_T_5 ? _GEN_27279 : rob_uop_13_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29714 = _next_will_commit_0_T_5 ? _GEN_27280 : rob_uop_14_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29715 = _next_will_commit_0_T_5 ? _GEN_27281 : rob_uop_15_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29716 = _next_will_commit_0_T_5 ? _GEN_27282 : rob_uop_16_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29717 = _next_will_commit_0_T_5 ? _GEN_27283 : rob_uop_17_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29718 = _next_will_commit_0_T_5 ? _GEN_27284 : rob_uop_18_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29719 = _next_will_commit_0_T_5 ? _GEN_27285 : rob_uop_19_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29720 = _next_will_commit_0_T_5 ? _GEN_27286 : rob_uop_20_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29721 = _next_will_commit_0_T_5 ? _GEN_27287 : rob_uop_21_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29722 = _next_will_commit_0_T_5 ? _GEN_27288 : rob_uop_22_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29723 = _next_will_commit_0_T_5 ? _GEN_27289 : rob_uop_23_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29724 = _next_will_commit_0_T_5 ? _GEN_27290 : rob_uop_24_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29725 = _next_will_commit_0_T_5 ? _GEN_27291 : rob_uop_25_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29726 = _next_will_commit_0_T_5 ? _GEN_27292 : rob_uop_26_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29727 = _next_will_commit_0_T_5 ? _GEN_27293 : rob_uop_27_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29728 = _next_will_commit_0_T_5 ? _GEN_27294 : rob_uop_28_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29729 = _next_will_commit_0_T_5 ? _GEN_27295 : rob_uop_29_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29730 = _next_will_commit_0_T_5 ? _GEN_27296 : rob_uop_30_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29731 = _next_will_commit_0_T_5 ? _GEN_27297 : rob_uop_31_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29732 = _next_will_commit_0_T_5 ? _GEN_27298 : rob_uop_32_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29733 = _next_will_commit_0_T_5 ? _GEN_27299 : rob_uop_33_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29734 = _next_will_commit_0_T_5 ? _GEN_27300 : rob_uop_34_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29735 = _next_will_commit_0_T_5 ? _GEN_27301 : rob_uop_35_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29736 = _next_will_commit_0_T_5 ? _GEN_27302 : rob_uop_36_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29737 = _next_will_commit_0_T_5 ? _GEN_27303 : rob_uop_37_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29738 = _next_will_commit_0_T_5 ? _GEN_27304 : rob_uop_38_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29739 = _next_will_commit_0_T_5 ? _GEN_27305 : rob_uop_39_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29740 = _next_will_commit_0_T_5 ? _GEN_27306 : rob_uop_40_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29741 = _next_will_commit_0_T_5 ? _GEN_27307 : rob_uop_41_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29742 = _next_will_commit_0_T_5 ? _GEN_27308 : rob_uop_42_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29743 = _next_will_commit_0_T_5 ? _GEN_27309 : rob_uop_43_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29744 = _next_will_commit_0_T_5 ? _GEN_27310 : rob_uop_44_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29745 = _next_will_commit_0_T_5 ? _GEN_27311 : rob_uop_45_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29746 = _next_will_commit_0_T_5 ? _GEN_27312 : rob_uop_46_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29747 = _next_will_commit_0_T_5 ? _GEN_27313 : rob_uop_47_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29748 = _next_will_commit_0_T_5 ? _GEN_27314 : rob_uop_48_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29749 = _next_will_commit_0_T_5 ? _GEN_27315 : rob_uop_49_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29750 = _next_will_commit_0_T_5 ? _GEN_27316 : rob_uop_50_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29751 = _next_will_commit_0_T_5 ? _GEN_27317 : rob_uop_51_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29752 = _next_will_commit_0_T_5 ? _GEN_27318 : rob_uop_52_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29753 = _next_will_commit_0_T_5 ? _GEN_27319 : rob_uop_53_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29754 = _next_will_commit_0_T_5 ? _GEN_27320 : rob_uop_54_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29755 = _next_will_commit_0_T_5 ? _GEN_27321 : rob_uop_55_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29756 = _next_will_commit_0_T_5 ? _GEN_27322 : rob_uop_56_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29757 = _next_will_commit_0_T_5 ? _GEN_27323 : rob_uop_57_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29758 = _next_will_commit_0_T_5 ? _GEN_27324 : rob_uop_58_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29759 = _next_will_commit_0_T_5 ? _GEN_27325 : rob_uop_59_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29760 = _next_will_commit_0_T_5 ? _GEN_27326 : rob_uop_60_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29761 = _next_will_commit_0_T_5 ? _GEN_27327 : rob_uop_61_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29762 = _next_will_commit_0_T_5 ? _GEN_27328 : rob_uop_62_src1_value; // @[rob.scala 123:38 82:26]
  wire [63:0] _GEN_29763 = _next_will_commit_0_T_5 ? _GEN_27329 : rob_uop_63_src1_value; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30020 = _next_will_commit_0_T_5 ? _GEN_27586 : rob_uop_0_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30021 = _next_will_commit_0_T_5 ? _GEN_27587 : rob_uop_1_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30022 = _next_will_commit_0_T_5 ? _GEN_27588 : rob_uop_2_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30023 = _next_will_commit_0_T_5 ? _GEN_27589 : rob_uop_3_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30024 = _next_will_commit_0_T_5 ? _GEN_27590 : rob_uop_4_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30025 = _next_will_commit_0_T_5 ? _GEN_27591 : rob_uop_5_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30026 = _next_will_commit_0_T_5 ? _GEN_27592 : rob_uop_6_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30027 = _next_will_commit_0_T_5 ? _GEN_27593 : rob_uop_7_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30028 = _next_will_commit_0_T_5 ? _GEN_27594 : rob_uop_8_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30029 = _next_will_commit_0_T_5 ? _GEN_27595 : rob_uop_9_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30030 = _next_will_commit_0_T_5 ? _GEN_27596 : rob_uop_10_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30031 = _next_will_commit_0_T_5 ? _GEN_27597 : rob_uop_11_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30032 = _next_will_commit_0_T_5 ? _GEN_27598 : rob_uop_12_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30033 = _next_will_commit_0_T_5 ? _GEN_27599 : rob_uop_13_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30034 = _next_will_commit_0_T_5 ? _GEN_27600 : rob_uop_14_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30035 = _next_will_commit_0_T_5 ? _GEN_27601 : rob_uop_15_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30036 = _next_will_commit_0_T_5 ? _GEN_27602 : rob_uop_16_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30037 = _next_will_commit_0_T_5 ? _GEN_27603 : rob_uop_17_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30038 = _next_will_commit_0_T_5 ? _GEN_27604 : rob_uop_18_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30039 = _next_will_commit_0_T_5 ? _GEN_27605 : rob_uop_19_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30040 = _next_will_commit_0_T_5 ? _GEN_27606 : rob_uop_20_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30041 = _next_will_commit_0_T_5 ? _GEN_27607 : rob_uop_21_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30042 = _next_will_commit_0_T_5 ? _GEN_27608 : rob_uop_22_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30043 = _next_will_commit_0_T_5 ? _GEN_27609 : rob_uop_23_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30044 = _next_will_commit_0_T_5 ? _GEN_27610 : rob_uop_24_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30045 = _next_will_commit_0_T_5 ? _GEN_27611 : rob_uop_25_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30046 = _next_will_commit_0_T_5 ? _GEN_27612 : rob_uop_26_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30047 = _next_will_commit_0_T_5 ? _GEN_27613 : rob_uop_27_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30048 = _next_will_commit_0_T_5 ? _GEN_27614 : rob_uop_28_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30049 = _next_will_commit_0_T_5 ? _GEN_27615 : rob_uop_29_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30050 = _next_will_commit_0_T_5 ? _GEN_27616 : rob_uop_30_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30051 = _next_will_commit_0_T_5 ? _GEN_27617 : rob_uop_31_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30052 = _next_will_commit_0_T_5 ? _GEN_27618 : rob_uop_32_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30053 = _next_will_commit_0_T_5 ? _GEN_27619 : rob_uop_33_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30054 = _next_will_commit_0_T_5 ? _GEN_27620 : rob_uop_34_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30055 = _next_will_commit_0_T_5 ? _GEN_27621 : rob_uop_35_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30056 = _next_will_commit_0_T_5 ? _GEN_27622 : rob_uop_36_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30057 = _next_will_commit_0_T_5 ? _GEN_27623 : rob_uop_37_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30058 = _next_will_commit_0_T_5 ? _GEN_27624 : rob_uop_38_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30059 = _next_will_commit_0_T_5 ? _GEN_27625 : rob_uop_39_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30060 = _next_will_commit_0_T_5 ? _GEN_27626 : rob_uop_40_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30061 = _next_will_commit_0_T_5 ? _GEN_27627 : rob_uop_41_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30062 = _next_will_commit_0_T_5 ? _GEN_27628 : rob_uop_42_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30063 = _next_will_commit_0_T_5 ? _GEN_27629 : rob_uop_43_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30064 = _next_will_commit_0_T_5 ? _GEN_27630 : rob_uop_44_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30065 = _next_will_commit_0_T_5 ? _GEN_27631 : rob_uop_45_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30066 = _next_will_commit_0_T_5 ? _GEN_27632 : rob_uop_46_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30067 = _next_will_commit_0_T_5 ? _GEN_27633 : rob_uop_47_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30068 = _next_will_commit_0_T_5 ? _GEN_27634 : rob_uop_48_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30069 = _next_will_commit_0_T_5 ? _GEN_27635 : rob_uop_49_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30070 = _next_will_commit_0_T_5 ? _GEN_27636 : rob_uop_50_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30071 = _next_will_commit_0_T_5 ? _GEN_27637 : rob_uop_51_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30072 = _next_will_commit_0_T_5 ? _GEN_27638 : rob_uop_52_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30073 = _next_will_commit_0_T_5 ? _GEN_27639 : rob_uop_53_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30074 = _next_will_commit_0_T_5 ? _GEN_27640 : rob_uop_54_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30075 = _next_will_commit_0_T_5 ? _GEN_27641 : rob_uop_55_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30076 = _next_will_commit_0_T_5 ? _GEN_27642 : rob_uop_56_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30077 = _next_will_commit_0_T_5 ? _GEN_27643 : rob_uop_57_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30078 = _next_will_commit_0_T_5 ? _GEN_27644 : rob_uop_58_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30079 = _next_will_commit_0_T_5 ? _GEN_27645 : rob_uop_59_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30080 = _next_will_commit_0_T_5 ? _GEN_27646 : rob_uop_60_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30081 = _next_will_commit_0_T_5 ? _GEN_27647 : rob_uop_61_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30082 = _next_will_commit_0_T_5 ? _GEN_27648 : rob_uop_62_alu_sel; // @[rob.scala 123:38 82:26]
  wire [4:0] _GEN_30083 = _next_will_commit_0_T_5 ? _GEN_27649 : rob_uop_63_alu_sel; // @[rob.scala 123:38 82:26]
  wire  _GEN_30212 = _next_will_commit_0_T_5 ? _GEN_28163 : rob_valid_0; // @[rob.scala 123:38 81:28]
  wire  _GEN_30213 = _next_will_commit_0_T_5 ? _GEN_28164 : rob_valid_1; // @[rob.scala 123:38 81:28]
  wire  _GEN_30214 = _next_will_commit_0_T_5 ? _GEN_28165 : rob_valid_2; // @[rob.scala 123:38 81:28]
  wire  _GEN_30215 = _next_will_commit_0_T_5 ? _GEN_28166 : rob_valid_3; // @[rob.scala 123:38 81:28]
  wire  _GEN_30216 = _next_will_commit_0_T_5 ? _GEN_28167 : rob_valid_4; // @[rob.scala 123:38 81:28]
  wire  _GEN_30217 = _next_will_commit_0_T_5 ? _GEN_28168 : rob_valid_5; // @[rob.scala 123:38 81:28]
  wire  _GEN_30218 = _next_will_commit_0_T_5 ? _GEN_28169 : rob_valid_6; // @[rob.scala 123:38 81:28]
  wire  _GEN_30219 = _next_will_commit_0_T_5 ? _GEN_28170 : rob_valid_7; // @[rob.scala 123:38 81:28]
  wire  _GEN_30220 = _next_will_commit_0_T_5 ? _GEN_28171 : rob_valid_8; // @[rob.scala 123:38 81:28]
  wire  _GEN_30221 = _next_will_commit_0_T_5 ? _GEN_28172 : rob_valid_9; // @[rob.scala 123:38 81:28]
  wire  _GEN_30222 = _next_will_commit_0_T_5 ? _GEN_28173 : rob_valid_10; // @[rob.scala 123:38 81:28]
  wire  _GEN_30223 = _next_will_commit_0_T_5 ? _GEN_28174 : rob_valid_11; // @[rob.scala 123:38 81:28]
  wire  _GEN_30224 = _next_will_commit_0_T_5 ? _GEN_28175 : rob_valid_12; // @[rob.scala 123:38 81:28]
  wire  _GEN_30225 = _next_will_commit_0_T_5 ? _GEN_28176 : rob_valid_13; // @[rob.scala 123:38 81:28]
  wire  _GEN_30226 = _next_will_commit_0_T_5 ? _GEN_28177 : rob_valid_14; // @[rob.scala 123:38 81:28]
  wire  _GEN_30227 = _next_will_commit_0_T_5 ? _GEN_28178 : rob_valid_15; // @[rob.scala 123:38 81:28]
  wire  _GEN_30228 = _next_will_commit_0_T_5 ? _GEN_28179 : rob_valid_16; // @[rob.scala 123:38 81:28]
  wire  _GEN_30229 = _next_will_commit_0_T_5 ? _GEN_28180 : rob_valid_17; // @[rob.scala 123:38 81:28]
  wire  _GEN_30230 = _next_will_commit_0_T_5 ? _GEN_28181 : rob_valid_18; // @[rob.scala 123:38 81:28]
  wire  _GEN_30231 = _next_will_commit_0_T_5 ? _GEN_28182 : rob_valid_19; // @[rob.scala 123:38 81:28]
  wire  _GEN_30232 = _next_will_commit_0_T_5 ? _GEN_28183 : rob_valid_20; // @[rob.scala 123:38 81:28]
  wire  _GEN_30233 = _next_will_commit_0_T_5 ? _GEN_28184 : rob_valid_21; // @[rob.scala 123:38 81:28]
  wire  _GEN_30234 = _next_will_commit_0_T_5 ? _GEN_28185 : rob_valid_22; // @[rob.scala 123:38 81:28]
  wire  _GEN_30235 = _next_will_commit_0_T_5 ? _GEN_28186 : rob_valid_23; // @[rob.scala 123:38 81:28]
  wire  _GEN_30236 = _next_will_commit_0_T_5 ? _GEN_28187 : rob_valid_24; // @[rob.scala 123:38 81:28]
  wire  _GEN_30237 = _next_will_commit_0_T_5 ? _GEN_28188 : rob_valid_25; // @[rob.scala 123:38 81:28]
  wire  _GEN_30238 = _next_will_commit_0_T_5 ? _GEN_28189 : rob_valid_26; // @[rob.scala 123:38 81:28]
  wire  _GEN_30239 = _next_will_commit_0_T_5 ? _GEN_28190 : rob_valid_27; // @[rob.scala 123:38 81:28]
  wire  _GEN_30240 = _next_will_commit_0_T_5 ? _GEN_28191 : rob_valid_28; // @[rob.scala 123:38 81:28]
  wire  _GEN_30241 = _next_will_commit_0_T_5 ? _GEN_28192 : rob_valid_29; // @[rob.scala 123:38 81:28]
  wire  _GEN_30242 = _next_will_commit_0_T_5 ? _GEN_28193 : rob_valid_30; // @[rob.scala 123:38 81:28]
  wire  _GEN_30243 = _next_will_commit_0_T_5 ? _GEN_28194 : rob_valid_31; // @[rob.scala 123:38 81:28]
  wire  _GEN_30244 = _next_will_commit_0_T_5 ? _GEN_28195 : rob_valid_32; // @[rob.scala 123:38 81:28]
  wire  _GEN_30245 = _next_will_commit_0_T_5 ? _GEN_28196 : rob_valid_33; // @[rob.scala 123:38 81:28]
  wire  _GEN_30246 = _next_will_commit_0_T_5 ? _GEN_28197 : rob_valid_34; // @[rob.scala 123:38 81:28]
  wire  _GEN_30247 = _next_will_commit_0_T_5 ? _GEN_28198 : rob_valid_35; // @[rob.scala 123:38 81:28]
  wire  _GEN_30248 = _next_will_commit_0_T_5 ? _GEN_28199 : rob_valid_36; // @[rob.scala 123:38 81:28]
  wire  _GEN_30249 = _next_will_commit_0_T_5 ? _GEN_28200 : rob_valid_37; // @[rob.scala 123:38 81:28]
  wire  _GEN_30250 = _next_will_commit_0_T_5 ? _GEN_28201 : rob_valid_38; // @[rob.scala 123:38 81:28]
  wire  _GEN_30251 = _next_will_commit_0_T_5 ? _GEN_28202 : rob_valid_39; // @[rob.scala 123:38 81:28]
  wire  _GEN_30252 = _next_will_commit_0_T_5 ? _GEN_28203 : rob_valid_40; // @[rob.scala 123:38 81:28]
  wire  _GEN_30253 = _next_will_commit_0_T_5 ? _GEN_28204 : rob_valid_41; // @[rob.scala 123:38 81:28]
  wire  _GEN_30254 = _next_will_commit_0_T_5 ? _GEN_28205 : rob_valid_42; // @[rob.scala 123:38 81:28]
  wire  _GEN_30255 = _next_will_commit_0_T_5 ? _GEN_28206 : rob_valid_43; // @[rob.scala 123:38 81:28]
  wire  _GEN_30256 = _next_will_commit_0_T_5 ? _GEN_28207 : rob_valid_44; // @[rob.scala 123:38 81:28]
  wire  _GEN_30257 = _next_will_commit_0_T_5 ? _GEN_28208 : rob_valid_45; // @[rob.scala 123:38 81:28]
  wire  _GEN_30258 = _next_will_commit_0_T_5 ? _GEN_28209 : rob_valid_46; // @[rob.scala 123:38 81:28]
  wire  _GEN_30259 = _next_will_commit_0_T_5 ? _GEN_28210 : rob_valid_47; // @[rob.scala 123:38 81:28]
  wire  _GEN_30260 = _next_will_commit_0_T_5 ? _GEN_28211 : rob_valid_48; // @[rob.scala 123:38 81:28]
  wire  _GEN_30261 = _next_will_commit_0_T_5 ? _GEN_28212 : rob_valid_49; // @[rob.scala 123:38 81:28]
  wire  _GEN_30262 = _next_will_commit_0_T_5 ? _GEN_28213 : rob_valid_50; // @[rob.scala 123:38 81:28]
  wire  _GEN_30263 = _next_will_commit_0_T_5 ? _GEN_28214 : rob_valid_51; // @[rob.scala 123:38 81:28]
  wire  _GEN_30264 = _next_will_commit_0_T_5 ? _GEN_28215 : rob_valid_52; // @[rob.scala 123:38 81:28]
  wire  _GEN_30265 = _next_will_commit_0_T_5 ? _GEN_28216 : rob_valid_53; // @[rob.scala 123:38 81:28]
  wire  _GEN_30266 = _next_will_commit_0_T_5 ? _GEN_28217 : rob_valid_54; // @[rob.scala 123:38 81:28]
  wire  _GEN_30267 = _next_will_commit_0_T_5 ? _GEN_28218 : rob_valid_55; // @[rob.scala 123:38 81:28]
  wire  _GEN_30268 = _next_will_commit_0_T_5 ? _GEN_28219 : rob_valid_56; // @[rob.scala 123:38 81:28]
  wire  _GEN_30269 = _next_will_commit_0_T_5 ? _GEN_28220 : rob_valid_57; // @[rob.scala 123:38 81:28]
  wire  _GEN_30270 = _next_will_commit_0_T_5 ? _GEN_28221 : rob_valid_58; // @[rob.scala 123:38 81:28]
  wire  _GEN_30271 = _next_will_commit_0_T_5 ? _GEN_28222 : rob_valid_59; // @[rob.scala 123:38 81:28]
  wire  _GEN_30272 = _next_will_commit_0_T_5 ? _GEN_28223 : rob_valid_60; // @[rob.scala 123:38 81:28]
  wire  _GEN_30273 = _next_will_commit_0_T_5 ? _GEN_28224 : rob_valid_61; // @[rob.scala 123:38 81:28]
  wire  _GEN_30274 = _next_will_commit_0_T_5 ? _GEN_28225 : rob_valid_62; // @[rob.scala 123:38 81:28]
  wire  _GEN_30275 = _next_will_commit_0_T_5 ? _GEN_28226 : rob_valid_63; // @[rob.scala 123:38 81:28]
  wire  _GEN_30276 = _next_will_commit_0_T_5 ? _GEN_27842 : rob_done_0; // @[rob.scala 123:38 84:27]
  wire  _GEN_30277 = _next_will_commit_0_T_5 ? _GEN_27843 : rob_done_1; // @[rob.scala 123:38 84:27]
  wire  _GEN_30278 = _next_will_commit_0_T_5 ? _GEN_27844 : rob_done_2; // @[rob.scala 123:38 84:27]
  wire  _GEN_30279 = _next_will_commit_0_T_5 ? _GEN_27845 : rob_done_3; // @[rob.scala 123:38 84:27]
  wire  _GEN_30280 = _next_will_commit_0_T_5 ? _GEN_27846 : rob_done_4; // @[rob.scala 123:38 84:27]
  wire  _GEN_30281 = _next_will_commit_0_T_5 ? _GEN_27847 : rob_done_5; // @[rob.scala 123:38 84:27]
  wire  _GEN_30282 = _next_will_commit_0_T_5 ? _GEN_27848 : rob_done_6; // @[rob.scala 123:38 84:27]
  wire  _GEN_30283 = _next_will_commit_0_T_5 ? _GEN_27849 : rob_done_7; // @[rob.scala 123:38 84:27]
  wire  _GEN_30284 = _next_will_commit_0_T_5 ? _GEN_27850 : rob_done_8; // @[rob.scala 123:38 84:27]
  wire  _GEN_30285 = _next_will_commit_0_T_5 ? _GEN_27851 : rob_done_9; // @[rob.scala 123:38 84:27]
  wire  _GEN_30286 = _next_will_commit_0_T_5 ? _GEN_27852 : rob_done_10; // @[rob.scala 123:38 84:27]
  wire  _GEN_30287 = _next_will_commit_0_T_5 ? _GEN_27853 : rob_done_11; // @[rob.scala 123:38 84:27]
  wire  _GEN_30288 = _next_will_commit_0_T_5 ? _GEN_27854 : rob_done_12; // @[rob.scala 123:38 84:27]
  wire  _GEN_30289 = _next_will_commit_0_T_5 ? _GEN_27855 : rob_done_13; // @[rob.scala 123:38 84:27]
  wire  _GEN_30290 = _next_will_commit_0_T_5 ? _GEN_27856 : rob_done_14; // @[rob.scala 123:38 84:27]
  wire  _GEN_30291 = _next_will_commit_0_T_5 ? _GEN_27857 : rob_done_15; // @[rob.scala 123:38 84:27]
  wire  _GEN_30292 = _next_will_commit_0_T_5 ? _GEN_27858 : rob_done_16; // @[rob.scala 123:38 84:27]
  wire  _GEN_30293 = _next_will_commit_0_T_5 ? _GEN_27859 : rob_done_17; // @[rob.scala 123:38 84:27]
  wire  _GEN_30294 = _next_will_commit_0_T_5 ? _GEN_27860 : rob_done_18; // @[rob.scala 123:38 84:27]
  wire  _GEN_30295 = _next_will_commit_0_T_5 ? _GEN_27861 : rob_done_19; // @[rob.scala 123:38 84:27]
  wire  _GEN_30296 = _next_will_commit_0_T_5 ? _GEN_27862 : rob_done_20; // @[rob.scala 123:38 84:27]
  wire  _GEN_30297 = _next_will_commit_0_T_5 ? _GEN_27863 : rob_done_21; // @[rob.scala 123:38 84:27]
  wire  _GEN_30298 = _next_will_commit_0_T_5 ? _GEN_27864 : rob_done_22; // @[rob.scala 123:38 84:27]
  wire  _GEN_30299 = _next_will_commit_0_T_5 ? _GEN_27865 : rob_done_23; // @[rob.scala 123:38 84:27]
  wire  _GEN_30300 = _next_will_commit_0_T_5 ? _GEN_27866 : rob_done_24; // @[rob.scala 123:38 84:27]
  wire  _GEN_30301 = _next_will_commit_0_T_5 ? _GEN_27867 : rob_done_25; // @[rob.scala 123:38 84:27]
  wire  _GEN_30302 = _next_will_commit_0_T_5 ? _GEN_27868 : rob_done_26; // @[rob.scala 123:38 84:27]
  wire  _GEN_30303 = _next_will_commit_0_T_5 ? _GEN_27869 : rob_done_27; // @[rob.scala 123:38 84:27]
  wire  _GEN_30304 = _next_will_commit_0_T_5 ? _GEN_27870 : rob_done_28; // @[rob.scala 123:38 84:27]
  wire  _GEN_30305 = _next_will_commit_0_T_5 ? _GEN_27871 : rob_done_29; // @[rob.scala 123:38 84:27]
  wire  _GEN_30306 = _next_will_commit_0_T_5 ? _GEN_27872 : rob_done_30; // @[rob.scala 123:38 84:27]
  wire  _GEN_30307 = _next_will_commit_0_T_5 ? _GEN_27873 : rob_done_31; // @[rob.scala 123:38 84:27]
  wire  _GEN_30308 = _next_will_commit_0_T_5 ? _GEN_27874 : rob_done_32; // @[rob.scala 123:38 84:27]
  wire  _GEN_30309 = _next_will_commit_0_T_5 ? _GEN_27875 : rob_done_33; // @[rob.scala 123:38 84:27]
  wire  _GEN_30310 = _next_will_commit_0_T_5 ? _GEN_27876 : rob_done_34; // @[rob.scala 123:38 84:27]
  wire  _GEN_30311 = _next_will_commit_0_T_5 ? _GEN_27877 : rob_done_35; // @[rob.scala 123:38 84:27]
  wire  _GEN_30312 = _next_will_commit_0_T_5 ? _GEN_27878 : rob_done_36; // @[rob.scala 123:38 84:27]
  wire  _GEN_30313 = _next_will_commit_0_T_5 ? _GEN_27879 : rob_done_37; // @[rob.scala 123:38 84:27]
  wire  _GEN_30314 = _next_will_commit_0_T_5 ? _GEN_27880 : rob_done_38; // @[rob.scala 123:38 84:27]
  wire  _GEN_30315 = _next_will_commit_0_T_5 ? _GEN_27881 : rob_done_39; // @[rob.scala 123:38 84:27]
  wire  _GEN_30316 = _next_will_commit_0_T_5 ? _GEN_27882 : rob_done_40; // @[rob.scala 123:38 84:27]
  wire  _GEN_30317 = _next_will_commit_0_T_5 ? _GEN_27883 : rob_done_41; // @[rob.scala 123:38 84:27]
  wire  _GEN_30318 = _next_will_commit_0_T_5 ? _GEN_27884 : rob_done_42; // @[rob.scala 123:38 84:27]
  wire  _GEN_30319 = _next_will_commit_0_T_5 ? _GEN_27885 : rob_done_43; // @[rob.scala 123:38 84:27]
  wire  _GEN_30320 = _next_will_commit_0_T_5 ? _GEN_27886 : rob_done_44; // @[rob.scala 123:38 84:27]
  wire  _GEN_30321 = _next_will_commit_0_T_5 ? _GEN_27887 : rob_done_45; // @[rob.scala 123:38 84:27]
  wire  _GEN_30322 = _next_will_commit_0_T_5 ? _GEN_27888 : rob_done_46; // @[rob.scala 123:38 84:27]
  wire  _GEN_30323 = _next_will_commit_0_T_5 ? _GEN_27889 : rob_done_47; // @[rob.scala 123:38 84:27]
  wire  _GEN_30324 = _next_will_commit_0_T_5 ? _GEN_27890 : rob_done_48; // @[rob.scala 123:38 84:27]
  wire  _GEN_30325 = _next_will_commit_0_T_5 ? _GEN_27891 : rob_done_49; // @[rob.scala 123:38 84:27]
  wire  _GEN_30326 = _next_will_commit_0_T_5 ? _GEN_27892 : rob_done_50; // @[rob.scala 123:38 84:27]
  wire  _GEN_30327 = _next_will_commit_0_T_5 ? _GEN_27893 : rob_done_51; // @[rob.scala 123:38 84:27]
  wire  _GEN_30328 = _next_will_commit_0_T_5 ? _GEN_27894 : rob_done_52; // @[rob.scala 123:38 84:27]
  wire  _GEN_30329 = _next_will_commit_0_T_5 ? _GEN_27895 : rob_done_53; // @[rob.scala 123:38 84:27]
  wire  _GEN_30330 = _next_will_commit_0_T_5 ? _GEN_27896 : rob_done_54; // @[rob.scala 123:38 84:27]
  wire  _GEN_30331 = _next_will_commit_0_T_5 ? _GEN_27897 : rob_done_55; // @[rob.scala 123:38 84:27]
  wire  _GEN_30332 = _next_will_commit_0_T_5 ? _GEN_27898 : rob_done_56; // @[rob.scala 123:38 84:27]
  wire  _GEN_30333 = _next_will_commit_0_T_5 ? _GEN_27899 : rob_done_57; // @[rob.scala 123:38 84:27]
  wire  _GEN_30334 = _next_will_commit_0_T_5 ? _GEN_27900 : rob_done_58; // @[rob.scala 123:38 84:27]
  wire  _GEN_30335 = _next_will_commit_0_T_5 ? _GEN_27901 : rob_done_59; // @[rob.scala 123:38 84:27]
  wire  _GEN_30336 = _next_will_commit_0_T_5 ? _GEN_27902 : rob_done_60; // @[rob.scala 123:38 84:27]
  wire  _GEN_30337 = _next_will_commit_0_T_5 ? _GEN_27903 : rob_done_61; // @[rob.scala 123:38 84:27]
  wire  _GEN_30338 = _next_will_commit_0_T_5 ? _GEN_27904 : rob_done_62; // @[rob.scala 123:38 84:27]
  wire  _GEN_30339 = _next_will_commit_0_T_5 ? _GEN_27905 : rob_done_63; // @[rob.scala 123:38 84:27]
  wire [6:0] _GEN_30405 = _next_will_commit_0_T_5 ? _GEN_28227 : commit_ptr; // @[rob.scala 123:38 46:29]
  wire  _GEN_30406 = _GEN_42065 | _GEN_30212; // @[rob.scala 167:{53,53}]
  wire  _GEN_30407 = _GEN_42066 | _GEN_30213; // @[rob.scala 167:{53,53}]
  wire  _GEN_30408 = _GEN_42067 | _GEN_30214; // @[rob.scala 167:{53,53}]
  wire  _GEN_30409 = _GEN_42068 | _GEN_30215; // @[rob.scala 167:{53,53}]
  wire  _GEN_30410 = _GEN_42069 | _GEN_30216; // @[rob.scala 167:{53,53}]
  wire  _GEN_30411 = _GEN_42070 | _GEN_30217; // @[rob.scala 167:{53,53}]
  wire  _GEN_30412 = _GEN_42071 | _GEN_30218; // @[rob.scala 167:{53,53}]
  wire  _GEN_30413 = _GEN_42072 | _GEN_30219; // @[rob.scala 167:{53,53}]
  wire  _GEN_30414 = _GEN_42073 | _GEN_30220; // @[rob.scala 167:{53,53}]
  wire  _GEN_30415 = _GEN_42074 | _GEN_30221; // @[rob.scala 167:{53,53}]
  wire  _GEN_30416 = _GEN_42075 | _GEN_30222; // @[rob.scala 167:{53,53}]
  wire  _GEN_30417 = _GEN_42076 | _GEN_30223; // @[rob.scala 167:{53,53}]
  wire  _GEN_30418 = _GEN_42077 | _GEN_30224; // @[rob.scala 167:{53,53}]
  wire  _GEN_30419 = _GEN_42078 | _GEN_30225; // @[rob.scala 167:{53,53}]
  wire  _GEN_30420 = _GEN_42079 | _GEN_30226; // @[rob.scala 167:{53,53}]
  wire  _GEN_30421 = _GEN_42080 | _GEN_30227; // @[rob.scala 167:{53,53}]
  wire  _GEN_30422 = _GEN_42081 | _GEN_30228; // @[rob.scala 167:{53,53}]
  wire  _GEN_30423 = _GEN_42082 | _GEN_30229; // @[rob.scala 167:{53,53}]
  wire  _GEN_30424 = _GEN_42083 | _GEN_30230; // @[rob.scala 167:{53,53}]
  wire  _GEN_30425 = _GEN_42084 | _GEN_30231; // @[rob.scala 167:{53,53}]
  wire  _GEN_30426 = _GEN_42085 | _GEN_30232; // @[rob.scala 167:{53,53}]
  wire  _GEN_30427 = _GEN_42086 | _GEN_30233; // @[rob.scala 167:{53,53}]
  wire  _GEN_30428 = _GEN_42087 | _GEN_30234; // @[rob.scala 167:{53,53}]
  wire  _GEN_30429 = _GEN_42088 | _GEN_30235; // @[rob.scala 167:{53,53}]
  wire  _GEN_30430 = _GEN_42089 | _GEN_30236; // @[rob.scala 167:{53,53}]
  wire  _GEN_30431 = _GEN_42090 | _GEN_30237; // @[rob.scala 167:{53,53}]
  wire  _GEN_30432 = _GEN_42091 | _GEN_30238; // @[rob.scala 167:{53,53}]
  wire  _GEN_30433 = _GEN_42092 | _GEN_30239; // @[rob.scala 167:{53,53}]
  wire  _GEN_30434 = _GEN_42093 | _GEN_30240; // @[rob.scala 167:{53,53}]
  wire  _GEN_30435 = _GEN_42094 | _GEN_30241; // @[rob.scala 167:{53,53}]
  wire  _GEN_30436 = _GEN_42095 | _GEN_30242; // @[rob.scala 167:{53,53}]
  wire  _GEN_30437 = _GEN_42096 | _GEN_30243; // @[rob.scala 167:{53,53}]
  wire  _GEN_30438 = _GEN_42097 | _GEN_30244; // @[rob.scala 167:{53,53}]
  wire  _GEN_30439 = _GEN_42098 | _GEN_30245; // @[rob.scala 167:{53,53}]
  wire  _GEN_30440 = _GEN_42099 | _GEN_30246; // @[rob.scala 167:{53,53}]
  wire  _GEN_30441 = _GEN_42100 | _GEN_30247; // @[rob.scala 167:{53,53}]
  wire  _GEN_30442 = _GEN_42101 | _GEN_30248; // @[rob.scala 167:{53,53}]
  wire  _GEN_30443 = _GEN_42102 | _GEN_30249; // @[rob.scala 167:{53,53}]
  wire  _GEN_30444 = _GEN_42103 | _GEN_30250; // @[rob.scala 167:{53,53}]
  wire  _GEN_30445 = _GEN_42104 | _GEN_30251; // @[rob.scala 167:{53,53}]
  wire  _GEN_30446 = _GEN_42105 | _GEN_30252; // @[rob.scala 167:{53,53}]
  wire  _GEN_30447 = _GEN_42106 | _GEN_30253; // @[rob.scala 167:{53,53}]
  wire  _GEN_30448 = _GEN_42107 | _GEN_30254; // @[rob.scala 167:{53,53}]
  wire  _GEN_30449 = _GEN_42108 | _GEN_30255; // @[rob.scala 167:{53,53}]
  wire  _GEN_30450 = _GEN_42109 | _GEN_30256; // @[rob.scala 167:{53,53}]
  wire  _GEN_30451 = _GEN_42110 | _GEN_30257; // @[rob.scala 167:{53,53}]
  wire  _GEN_30452 = _GEN_42111 | _GEN_30258; // @[rob.scala 167:{53,53}]
  wire  _GEN_30453 = _GEN_42112 | _GEN_30259; // @[rob.scala 167:{53,53}]
  wire  _GEN_30454 = _GEN_42113 | _GEN_30260; // @[rob.scala 167:{53,53}]
  wire  _GEN_30455 = _GEN_42114 | _GEN_30261; // @[rob.scala 167:{53,53}]
  wire  _GEN_30456 = _GEN_42115 | _GEN_30262; // @[rob.scala 167:{53,53}]
  wire  _GEN_30457 = _GEN_42116 | _GEN_30263; // @[rob.scala 167:{53,53}]
  wire  _GEN_30458 = _GEN_42117 | _GEN_30264; // @[rob.scala 167:{53,53}]
  wire  _GEN_30459 = _GEN_42118 | _GEN_30265; // @[rob.scala 167:{53,53}]
  wire  _GEN_30460 = _GEN_42119 | _GEN_30266; // @[rob.scala 167:{53,53}]
  wire  _GEN_30461 = _GEN_42120 | _GEN_30267; // @[rob.scala 167:{53,53}]
  wire  _GEN_30462 = _GEN_42121 | _GEN_30268; // @[rob.scala 167:{53,53}]
  wire  _GEN_30463 = _GEN_42122 | _GEN_30269; // @[rob.scala 167:{53,53}]
  wire  _GEN_30464 = _GEN_42123 | _GEN_30270; // @[rob.scala 167:{53,53}]
  wire  _GEN_30465 = _GEN_42124 | _GEN_30271; // @[rob.scala 167:{53,53}]
  wire  _GEN_30466 = _GEN_42125 | _GEN_30272; // @[rob.scala 167:{53,53}]
  wire  _GEN_30467 = _GEN_42126 | _GEN_30273; // @[rob.scala 167:{53,53}]
  wire  _GEN_30468 = _GEN_42127 | _GEN_30274; // @[rob.scala 167:{53,53}]
  wire  _GEN_30469 = _GEN_42128 | _GEN_30275; // @[rob.scala 167:{53,53}]
  wire [31:0] _GEN_30534 = 6'h0 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28292; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30535 = 6'h1 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28293; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30536 = 6'h2 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28294; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30537 = 6'h3 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28295; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30538 = 6'h4 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28296; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30539 = 6'h5 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28297; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30540 = 6'h6 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28298; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30541 = 6'h7 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28299; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30542 = 6'h8 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28300; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30543 = 6'h9 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28301; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30544 = 6'ha == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28302; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30545 = 6'hb == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28303; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30546 = 6'hc == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28304; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30547 = 6'hd == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28305; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30548 = 6'he == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28306; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30549 = 6'hf == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28307; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30550 = 6'h10 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28308; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30551 = 6'h11 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28309; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30552 = 6'h12 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28310; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30553 = 6'h13 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28311; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30554 = 6'h14 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28312; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30555 = 6'h15 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28313; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30556 = 6'h16 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28314; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30557 = 6'h17 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28315; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30558 = 6'h18 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28316; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30559 = 6'h19 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28317; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30560 = 6'h1a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28318; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30561 = 6'h1b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28319; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30562 = 6'h1c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28320; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30563 = 6'h1d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28321; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30564 = 6'h1e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28322; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30565 = 6'h1f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28323; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30566 = 6'h20 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28324; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30567 = 6'h21 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28325; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30568 = 6'h22 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28326; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30569 = 6'h23 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28327; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30570 = 6'h24 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28328; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30571 = 6'h25 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28329; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30572 = 6'h26 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28330; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30573 = 6'h27 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28331; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30574 = 6'h28 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28332; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30575 = 6'h29 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28333; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30576 = 6'h2a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28334; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30577 = 6'h2b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28335; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30578 = 6'h2c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28336; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30579 = 6'h2d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28337; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30580 = 6'h2e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28338; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30581 = 6'h2f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28339; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30582 = 6'h30 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28340; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30583 = 6'h31 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28341; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30584 = 6'h32 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28342; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30585 = 6'h33 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28343; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30586 = 6'h34 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28344; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30587 = 6'h35 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28345; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30588 = 6'h36 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28346; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30589 = 6'h37 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28347; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30590 = 6'h38 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28348; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30591 = 6'h39 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28349; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30592 = 6'h3a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28350; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30593 = 6'h3b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28351; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30594 = 6'h3c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28352; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30595 = 6'h3d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28353; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30596 = 6'h3e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28354; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30597 = 6'h3f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_pc : _GEN_28355; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30598 = 6'h0 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28356; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30599 = 6'h1 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28357; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30600 = 6'h2 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28358; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30601 = 6'h3 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28359; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30602 = 6'h4 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28360; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30603 = 6'h5 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28361; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30604 = 6'h6 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28362; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30605 = 6'h7 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28363; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30606 = 6'h8 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28364; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30607 = 6'h9 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28365; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30608 = 6'ha == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28366; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30609 = 6'hb == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28367; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30610 = 6'hc == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28368; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30611 = 6'hd == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28369; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30612 = 6'he == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28370; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30613 = 6'hf == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28371; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30614 = 6'h10 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28372; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30615 = 6'h11 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28373; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30616 = 6'h12 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28374; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30617 = 6'h13 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28375; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30618 = 6'h14 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28376; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30619 = 6'h15 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28377; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30620 = 6'h16 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28378; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30621 = 6'h17 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28379; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30622 = 6'h18 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28380; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30623 = 6'h19 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28381; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30624 = 6'h1a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28382; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30625 = 6'h1b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28383; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30626 = 6'h1c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28384; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30627 = 6'h1d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28385; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30628 = 6'h1e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28386; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30629 = 6'h1f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28387; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30630 = 6'h20 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28388; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30631 = 6'h21 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28389; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30632 = 6'h22 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28390; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30633 = 6'h23 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28391; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30634 = 6'h24 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28392; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30635 = 6'h25 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28393; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30636 = 6'h26 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28394; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30637 = 6'h27 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28395; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30638 = 6'h28 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28396; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30639 = 6'h29 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28397; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30640 = 6'h2a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28398; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30641 = 6'h2b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28399; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30642 = 6'h2c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28400; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30643 = 6'h2d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28401; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30644 = 6'h2e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28402; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30645 = 6'h2f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28403; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30646 = 6'h30 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28404; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30647 = 6'h31 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28405; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30648 = 6'h32 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28406; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30649 = 6'h33 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28407; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30650 = 6'h34 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28408; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30651 = 6'h35 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28409; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30652 = 6'h36 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28410; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30653 = 6'h37 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28411; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30654 = 6'h38 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28412; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30655 = 6'h39 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28413; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30656 = 6'h3a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28414; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30657 = 6'h3b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28415; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30658 = 6'h3c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28416; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30659 = 6'h3d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28417; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30660 = 6'h3e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28418; // @[rob.scala 168:{51,51}]
  wire [31:0] _GEN_30661 = 6'h3f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_inst : _GEN_28419; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30662 = 6'h0 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28420; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30663 = 6'h1 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28421; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30664 = 6'h2 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28422; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30665 = 6'h3 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28423; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30666 = 6'h4 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28424; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30667 = 6'h5 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28425; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30668 = 6'h6 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28426; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30669 = 6'h7 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28427; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30670 = 6'h8 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28428; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30671 = 6'h9 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28429; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30672 = 6'ha == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28430; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30673 = 6'hb == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28431; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30674 = 6'hc == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28432; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30675 = 6'hd == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28433; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30676 = 6'he == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28434; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30677 = 6'hf == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28435; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30678 = 6'h10 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28436
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30679 = 6'h11 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28437
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30680 = 6'h12 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28438
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30681 = 6'h13 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28439
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30682 = 6'h14 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28440
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30683 = 6'h15 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28441
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30684 = 6'h16 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28442
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30685 = 6'h17 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28443
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30686 = 6'h18 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28444
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30687 = 6'h19 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28445
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30688 = 6'h1a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28446
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30689 = 6'h1b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28447
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30690 = 6'h1c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28448
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30691 = 6'h1d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28449
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30692 = 6'h1e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28450
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30693 = 6'h1f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28451
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30694 = 6'h20 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28452
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30695 = 6'h21 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28453
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30696 = 6'h22 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28454
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30697 = 6'h23 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28455
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30698 = 6'h24 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28456
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30699 = 6'h25 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28457
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30700 = 6'h26 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28458
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30701 = 6'h27 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28459
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30702 = 6'h28 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28460
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30703 = 6'h29 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28461
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30704 = 6'h2a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28462
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30705 = 6'h2b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28463
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30706 = 6'h2c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28464
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30707 = 6'h2d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28465
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30708 = 6'h2e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28466
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30709 = 6'h2f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28467
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30710 = 6'h30 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28468
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30711 = 6'h31 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28469
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30712 = 6'h32 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28470
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30713 = 6'h33 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28471
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30714 = 6'h34 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28472
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30715 = 6'h35 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28473
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30716 = 6'h36 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28474
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30717 = 6'h37 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28475
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30718 = 6'h38 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28476
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30719 = 6'h39 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28477
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30720 = 6'h3a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28478
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30721 = 6'h3b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28479
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30722 = 6'h3c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28480
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30723 = 6'h3d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28481
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30724 = 6'h3e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28482
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_30725 = 6'h3f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_func_code : _GEN_28483
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31046 = 6'h0 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28804; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31047 = 6'h1 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28805; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31048 = 6'h2 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28806; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31049 = 6'h3 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28807; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31050 = 6'h4 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28808; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31051 = 6'h5 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28809; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31052 = 6'h6 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28810; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31053 = 6'h7 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28811; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31054 = 6'h8 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28812; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31055 = 6'h9 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28813; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31056 = 6'ha == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28814; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31057 = 6'hb == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28815; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31058 = 6'hc == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28816; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31059 = 6'hd == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28817; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31060 = 6'he == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28818; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31061 = 6'hf == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28819; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31062 = 6'h10 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28820; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31063 = 6'h11 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28821; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31064 = 6'h12 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28822; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31065 = 6'h13 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28823; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31066 = 6'h14 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28824; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31067 = 6'h15 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28825; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31068 = 6'h16 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28826; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31069 = 6'h17 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28827; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31070 = 6'h18 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28828; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31071 = 6'h19 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28829; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31072 = 6'h1a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28830; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31073 = 6'h1b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28831; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31074 = 6'h1c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28832; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31075 = 6'h1d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28833; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31076 = 6'h1e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28834; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31077 = 6'h1f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28835; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31078 = 6'h20 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28836; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31079 = 6'h21 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28837; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31080 = 6'h22 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28838; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31081 = 6'h23 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28839; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31082 = 6'h24 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28840; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31083 = 6'h25 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28841; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31084 = 6'h26 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28842; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31085 = 6'h27 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28843; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31086 = 6'h28 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28844; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31087 = 6'h29 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28845; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31088 = 6'h2a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28846; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31089 = 6'h2b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28847; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31090 = 6'h2c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28848; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31091 = 6'h2d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28849; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31092 = 6'h2e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28850; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31093 = 6'h2f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28851; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31094 = 6'h30 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28852; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31095 = 6'h31 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28853; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31096 = 6'h32 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28854; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31097 = 6'h33 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28855; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31098 = 6'h34 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28856; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31099 = 6'h35 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28857; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31100 = 6'h36 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28858; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31101 = 6'h37 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28859; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31102 = 6'h38 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28860; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31103 = 6'h39 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28861; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31104 = 6'h3a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28862; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31105 = 6'h3b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28863; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31106 = 6'h3c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28864; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31107 = 6'h3d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28865; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31108 = 6'h3e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28866; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31109 = 6'h3f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_phy_dst : _GEN_28867; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31110 = 6'h0 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28868; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31111 = 6'h1 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28869; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31112 = 6'h2 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28870; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31113 = 6'h3 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28871; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31114 = 6'h4 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28872; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31115 = 6'h5 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28873; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31116 = 6'h6 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28874; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31117 = 6'h7 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28875; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31118 = 6'h8 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28876; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31119 = 6'h9 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28877; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31120 = 6'ha == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28878; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31121 = 6'hb == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28879; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31122 = 6'hc == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28880; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31123 = 6'hd == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28881; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31124 = 6'he == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28882; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31125 = 6'hf == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28883; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31126 = 6'h10 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28884
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31127 = 6'h11 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28885
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31128 = 6'h12 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28886
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31129 = 6'h13 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28887
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31130 = 6'h14 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28888
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31131 = 6'h15 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28889
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31132 = 6'h16 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28890
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31133 = 6'h17 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28891
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31134 = 6'h18 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28892
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31135 = 6'h19 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28893
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31136 = 6'h1a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28894
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31137 = 6'h1b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28895
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31138 = 6'h1c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28896
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31139 = 6'h1d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28897
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31140 = 6'h1e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28898
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31141 = 6'h1f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28899
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31142 = 6'h20 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28900
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31143 = 6'h21 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28901
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31144 = 6'h22 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28902
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31145 = 6'h23 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28903
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31146 = 6'h24 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28904
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31147 = 6'h25 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28905
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31148 = 6'h26 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28906
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31149 = 6'h27 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28907
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31150 = 6'h28 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28908
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31151 = 6'h29 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28909
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31152 = 6'h2a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28910
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31153 = 6'h2b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28911
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31154 = 6'h2c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28912
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31155 = 6'h2d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28913
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31156 = 6'h2e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28914
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31157 = 6'h2f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28915
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31158 = 6'h30 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28916
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31159 = 6'h31 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28917
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31160 = 6'h32 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28918
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31161 = 6'h33 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28919
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31162 = 6'h34 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28920
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31163 = 6'h35 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28921
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31164 = 6'h36 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28922
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31165 = 6'h37 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28923
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31166 = 6'h38 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28924
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31167 = 6'h39 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28925
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31168 = 6'h3a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28926
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31169 = 6'h3b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28927
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31170 = 6'h3c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28928
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31171 = 6'h3d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28929
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31172 = 6'h3e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28930
    ; // @[rob.scala 168:{51,51}]
  wire [6:0] _GEN_31173 = 6'h3f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_stale_dst : _GEN_28931
    ; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31174 = 6'h0 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28932; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31175 = 6'h1 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28933; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31176 = 6'h2 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28934; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31177 = 6'h3 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28935; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31178 = 6'h4 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28936; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31179 = 6'h5 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28937; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31180 = 6'h6 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28938; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31181 = 6'h7 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28939; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31182 = 6'h8 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28940; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31183 = 6'h9 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28941; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31184 = 6'ha == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28942; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31185 = 6'hb == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28943; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31186 = 6'hc == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28944; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31187 = 6'hd == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28945; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31188 = 6'he == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28946; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31189 = 6'hf == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28947; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31190 = 6'h10 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28948; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31191 = 6'h11 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28949; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31192 = 6'h12 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28950; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31193 = 6'h13 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28951; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31194 = 6'h14 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28952; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31195 = 6'h15 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28953; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31196 = 6'h16 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28954; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31197 = 6'h17 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28955; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31198 = 6'h18 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28956; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31199 = 6'h19 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28957; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31200 = 6'h1a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28958; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31201 = 6'h1b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28959; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31202 = 6'h1c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28960; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31203 = 6'h1d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28961; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31204 = 6'h1e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28962; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31205 = 6'h1f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28963; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31206 = 6'h20 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28964; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31207 = 6'h21 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28965; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31208 = 6'h22 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28966; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31209 = 6'h23 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28967; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31210 = 6'h24 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28968; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31211 = 6'h25 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28969; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31212 = 6'h26 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28970; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31213 = 6'h27 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28971; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31214 = 6'h28 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28972; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31215 = 6'h29 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28973; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31216 = 6'h2a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28974; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31217 = 6'h2b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28975; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31218 = 6'h2c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28976; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31219 = 6'h2d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28977; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31220 = 6'h2e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28978; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31221 = 6'h2f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28979; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31222 = 6'h30 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28980; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31223 = 6'h31 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28981; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31224 = 6'h32 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28982; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31225 = 6'h33 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28983; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31226 = 6'h34 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28984; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31227 = 6'h35 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28985; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31228 = 6'h36 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28986; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31229 = 6'h37 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28987; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31230 = 6'h38 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28988; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31231 = 6'h39 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28989; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31232 = 6'h3a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28990; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31233 = 6'h3b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28991; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31234 = 6'h3c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28992; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31235 = 6'h3d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28993; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31236 = 6'h3e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28994; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_31237 = 6'h3f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_arch_dst : _GEN_28995; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31878 = 6'h0 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value : _GEN_29636
    ; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31879 = 6'h1 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value : _GEN_29637
    ; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31880 = 6'h2 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value : _GEN_29638
    ; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31881 = 6'h3 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value : _GEN_29639
    ; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31882 = 6'h4 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value : _GEN_29640
    ; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31883 = 6'h5 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value : _GEN_29641
    ; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31884 = 6'h6 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value : _GEN_29642
    ; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31885 = 6'h7 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value : _GEN_29643
    ; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31886 = 6'h8 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value : _GEN_29644
    ; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31887 = 6'h9 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value : _GEN_29645
    ; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31888 = 6'ha == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value : _GEN_29646
    ; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31889 = 6'hb == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value : _GEN_29647
    ; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31890 = 6'hc == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value : _GEN_29648
    ; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31891 = 6'hd == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value : _GEN_29649
    ; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31892 = 6'he == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value : _GEN_29650
    ; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31893 = 6'hf == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value : _GEN_29651
    ; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31894 = 6'h10 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29652; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31895 = 6'h11 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29653; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31896 = 6'h12 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29654; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31897 = 6'h13 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29655; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31898 = 6'h14 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29656; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31899 = 6'h15 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29657; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31900 = 6'h16 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29658; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31901 = 6'h17 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29659; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31902 = 6'h18 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29660; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31903 = 6'h19 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29661; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31904 = 6'h1a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29662; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31905 = 6'h1b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29663; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31906 = 6'h1c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29664; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31907 = 6'h1d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29665; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31908 = 6'h1e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29666; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31909 = 6'h1f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29667; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31910 = 6'h20 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29668; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31911 = 6'h21 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29669; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31912 = 6'h22 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29670; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31913 = 6'h23 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29671; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31914 = 6'h24 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29672; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31915 = 6'h25 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29673; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31916 = 6'h26 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29674; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31917 = 6'h27 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29675; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31918 = 6'h28 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29676; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31919 = 6'h29 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29677; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31920 = 6'h2a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29678; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31921 = 6'h2b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29679; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31922 = 6'h2c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29680; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31923 = 6'h2d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29681; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31924 = 6'h2e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29682; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31925 = 6'h2f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29683; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31926 = 6'h30 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29684; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31927 = 6'h31 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29685; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31928 = 6'h32 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29686; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31929 = 6'h33 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29687; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31930 = 6'h34 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29688; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31931 = 6'h35 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29689; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31932 = 6'h36 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29690; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31933 = 6'h37 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29691; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31934 = 6'h38 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29692; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31935 = 6'h39 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29693; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31936 = 6'h3a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29694; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31937 = 6'h3b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29695; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31938 = 6'h3c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29696; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31939 = 6'h3d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29697; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31940 = 6'h3e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29698; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31941 = 6'h3f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_dst_value :
    _GEN_29699; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31942 = 6'h0 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29700; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31943 = 6'h1 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29701; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31944 = 6'h2 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29702; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31945 = 6'h3 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29703; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31946 = 6'h4 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29704; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31947 = 6'h5 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29705; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31948 = 6'h6 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29706; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31949 = 6'h7 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29707; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31950 = 6'h8 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29708; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31951 = 6'h9 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29709; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31952 = 6'ha == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29710; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31953 = 6'hb == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29711; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31954 = 6'hc == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29712; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31955 = 6'hd == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29713; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31956 = 6'he == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29714; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31957 = 6'hf == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29715; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31958 = 6'h10 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29716; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31959 = 6'h11 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29717; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31960 = 6'h12 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29718; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31961 = 6'h13 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29719; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31962 = 6'h14 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29720; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31963 = 6'h15 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29721; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31964 = 6'h16 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29722; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31965 = 6'h17 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29723; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31966 = 6'h18 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29724; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31967 = 6'h19 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29725; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31968 = 6'h1a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29726; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31969 = 6'h1b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29727; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31970 = 6'h1c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29728; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31971 = 6'h1d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29729; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31972 = 6'h1e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29730; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31973 = 6'h1f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29731; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31974 = 6'h20 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29732; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31975 = 6'h21 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29733; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31976 = 6'h22 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29734; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31977 = 6'h23 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29735; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31978 = 6'h24 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29736; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31979 = 6'h25 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29737; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31980 = 6'h26 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29738; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31981 = 6'h27 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29739; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31982 = 6'h28 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29740; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31983 = 6'h29 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29741; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31984 = 6'h2a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29742; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31985 = 6'h2b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29743; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31986 = 6'h2c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29744; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31987 = 6'h2d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29745; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31988 = 6'h2e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29746; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31989 = 6'h2f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29747; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31990 = 6'h30 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29748; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31991 = 6'h31 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29749; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31992 = 6'h32 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29750; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31993 = 6'h33 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29751; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31994 = 6'h34 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29752; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31995 = 6'h35 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29753; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31996 = 6'h36 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29754; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31997 = 6'h37 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29755; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31998 = 6'h38 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29756; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_31999 = 6'h39 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29757; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_32000 = 6'h3a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29758; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_32001 = 6'h3b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29759; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_32002 = 6'h3c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29760; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_32003 = 6'h3d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29761; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_32004 = 6'h3e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29762; // @[rob.scala 168:{51,51}]
  wire [63:0] _GEN_32005 = 6'h3f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_src1_value :
    _GEN_29763; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32262 = 6'h0 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30020; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32263 = 6'h1 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30021; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32264 = 6'h2 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30022; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32265 = 6'h3 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30023; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32266 = 6'h4 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30024; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32267 = 6'h5 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30025; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32268 = 6'h6 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30026; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32269 = 6'h7 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30027; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32270 = 6'h8 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30028; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32271 = 6'h9 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30029; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32272 = 6'ha == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30030; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32273 = 6'hb == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30031; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32274 = 6'hc == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30032; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32275 = 6'hd == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30033; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32276 = 6'he == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30034; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32277 = 6'hf == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30035; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32278 = 6'h10 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30036; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32279 = 6'h11 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30037; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32280 = 6'h12 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30038; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32281 = 6'h13 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30039; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32282 = 6'h14 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30040; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32283 = 6'h15 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30041; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32284 = 6'h16 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30042; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32285 = 6'h17 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30043; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32286 = 6'h18 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30044; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32287 = 6'h19 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30045; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32288 = 6'h1a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30046; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32289 = 6'h1b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30047; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32290 = 6'h1c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30048; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32291 = 6'h1d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30049; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32292 = 6'h1e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30050; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32293 = 6'h1f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30051; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32294 = 6'h20 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30052; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32295 = 6'h21 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30053; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32296 = 6'h22 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30054; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32297 = 6'h23 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30055; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32298 = 6'h24 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30056; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32299 = 6'h25 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30057; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32300 = 6'h26 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30058; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32301 = 6'h27 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30059; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32302 = 6'h28 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30060; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32303 = 6'h29 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30061; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32304 = 6'h2a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30062; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32305 = 6'h2b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30063; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32306 = 6'h2c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30064; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32307 = 6'h2d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30065; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32308 = 6'h2e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30066; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32309 = 6'h2f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30067; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32310 = 6'h30 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30068; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32311 = 6'h31 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30069; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32312 = 6'h32 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30070; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32313 = 6'h33 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30071; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32314 = 6'h34 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30072; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32315 = 6'h35 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30073; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32316 = 6'h36 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30074; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32317 = 6'h37 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30075; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32318 = 6'h38 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30076; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32319 = 6'h39 == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30077; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32320 = 6'h3a == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30078; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32321 = 6'h3b == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30079; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32322 = 6'h3c == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30080; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32323 = 6'h3d == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30081; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32324 = 6'h3e == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30082; // @[rob.scala 168:{51,51}]
  wire [4:0] _GEN_32325 = 6'h3f == io_i_ex_res_packs_0_uop_rob_idx[5:0] ? io_i_ex_res_packs_0_uop_alu_sel : _GEN_30083; // @[rob.scala 168:{51,51}]
  wire  _GEN_32518 = _GEN_42065 | _GEN_30276; // @[rob.scala 170:{52,52}]
  wire  _GEN_32519 = _GEN_42066 | _GEN_30277; // @[rob.scala 170:{52,52}]
  wire  _GEN_32520 = _GEN_42067 | _GEN_30278; // @[rob.scala 170:{52,52}]
  wire  _GEN_32521 = _GEN_42068 | _GEN_30279; // @[rob.scala 170:{52,52}]
  wire  _GEN_32522 = _GEN_42069 | _GEN_30280; // @[rob.scala 170:{52,52}]
  wire  _GEN_32523 = _GEN_42070 | _GEN_30281; // @[rob.scala 170:{52,52}]
  wire  _GEN_32524 = _GEN_42071 | _GEN_30282; // @[rob.scala 170:{52,52}]
  wire  _GEN_32525 = _GEN_42072 | _GEN_30283; // @[rob.scala 170:{52,52}]
  wire  _GEN_32526 = _GEN_42073 | _GEN_30284; // @[rob.scala 170:{52,52}]
  wire  _GEN_32527 = _GEN_42074 | _GEN_30285; // @[rob.scala 170:{52,52}]
  wire  _GEN_32528 = _GEN_42075 | _GEN_30286; // @[rob.scala 170:{52,52}]
  wire  _GEN_32529 = _GEN_42076 | _GEN_30287; // @[rob.scala 170:{52,52}]
  wire  _GEN_32530 = _GEN_42077 | _GEN_30288; // @[rob.scala 170:{52,52}]
  wire  _GEN_32531 = _GEN_42078 | _GEN_30289; // @[rob.scala 170:{52,52}]
  wire  _GEN_32532 = _GEN_42079 | _GEN_30290; // @[rob.scala 170:{52,52}]
  wire  _GEN_32533 = _GEN_42080 | _GEN_30291; // @[rob.scala 170:{52,52}]
  wire  _GEN_32534 = _GEN_42081 | _GEN_30292; // @[rob.scala 170:{52,52}]
  wire  _GEN_32535 = _GEN_42082 | _GEN_30293; // @[rob.scala 170:{52,52}]
  wire  _GEN_32536 = _GEN_42083 | _GEN_30294; // @[rob.scala 170:{52,52}]
  wire  _GEN_32537 = _GEN_42084 | _GEN_30295; // @[rob.scala 170:{52,52}]
  wire  _GEN_32538 = _GEN_42085 | _GEN_30296; // @[rob.scala 170:{52,52}]
  wire  _GEN_32539 = _GEN_42086 | _GEN_30297; // @[rob.scala 170:{52,52}]
  wire  _GEN_32540 = _GEN_42087 | _GEN_30298; // @[rob.scala 170:{52,52}]
  wire  _GEN_32541 = _GEN_42088 | _GEN_30299; // @[rob.scala 170:{52,52}]
  wire  _GEN_32542 = _GEN_42089 | _GEN_30300; // @[rob.scala 170:{52,52}]
  wire  _GEN_32543 = _GEN_42090 | _GEN_30301; // @[rob.scala 170:{52,52}]
  wire  _GEN_32544 = _GEN_42091 | _GEN_30302; // @[rob.scala 170:{52,52}]
  wire  _GEN_32545 = _GEN_42092 | _GEN_30303; // @[rob.scala 170:{52,52}]
  wire  _GEN_32546 = _GEN_42093 | _GEN_30304; // @[rob.scala 170:{52,52}]
  wire  _GEN_32547 = _GEN_42094 | _GEN_30305; // @[rob.scala 170:{52,52}]
  wire  _GEN_32548 = _GEN_42095 | _GEN_30306; // @[rob.scala 170:{52,52}]
  wire  _GEN_32549 = _GEN_42096 | _GEN_30307; // @[rob.scala 170:{52,52}]
  wire  _GEN_32550 = _GEN_42097 | _GEN_30308; // @[rob.scala 170:{52,52}]
  wire  _GEN_32551 = _GEN_42098 | _GEN_30309; // @[rob.scala 170:{52,52}]
  wire  _GEN_32552 = _GEN_42099 | _GEN_30310; // @[rob.scala 170:{52,52}]
  wire  _GEN_32553 = _GEN_42100 | _GEN_30311; // @[rob.scala 170:{52,52}]
  wire  _GEN_32554 = _GEN_42101 | _GEN_30312; // @[rob.scala 170:{52,52}]
  wire  _GEN_32555 = _GEN_42102 | _GEN_30313; // @[rob.scala 170:{52,52}]
  wire  _GEN_32556 = _GEN_42103 | _GEN_30314; // @[rob.scala 170:{52,52}]
  wire  _GEN_32557 = _GEN_42104 | _GEN_30315; // @[rob.scala 170:{52,52}]
  wire  _GEN_32558 = _GEN_42105 | _GEN_30316; // @[rob.scala 170:{52,52}]
  wire  _GEN_32559 = _GEN_42106 | _GEN_30317; // @[rob.scala 170:{52,52}]
  wire  _GEN_32560 = _GEN_42107 | _GEN_30318; // @[rob.scala 170:{52,52}]
  wire  _GEN_32561 = _GEN_42108 | _GEN_30319; // @[rob.scala 170:{52,52}]
  wire  _GEN_32562 = _GEN_42109 | _GEN_30320; // @[rob.scala 170:{52,52}]
  wire  _GEN_32563 = _GEN_42110 | _GEN_30321; // @[rob.scala 170:{52,52}]
  wire  _GEN_32564 = _GEN_42111 | _GEN_30322; // @[rob.scala 170:{52,52}]
  wire  _GEN_32565 = _GEN_42112 | _GEN_30323; // @[rob.scala 170:{52,52}]
  wire  _GEN_32566 = _GEN_42113 | _GEN_30324; // @[rob.scala 170:{52,52}]
  wire  _GEN_32567 = _GEN_42114 | _GEN_30325; // @[rob.scala 170:{52,52}]
  wire  _GEN_32568 = _GEN_42115 | _GEN_30326; // @[rob.scala 170:{52,52}]
  wire  _GEN_32569 = _GEN_42116 | _GEN_30327; // @[rob.scala 170:{52,52}]
  wire  _GEN_32570 = _GEN_42117 | _GEN_30328; // @[rob.scala 170:{52,52}]
  wire  _GEN_32571 = _GEN_42118 | _GEN_30329; // @[rob.scala 170:{52,52}]
  wire  _GEN_32572 = _GEN_42119 | _GEN_30330; // @[rob.scala 170:{52,52}]
  wire  _GEN_32573 = _GEN_42120 | _GEN_30331; // @[rob.scala 170:{52,52}]
  wire  _GEN_32574 = _GEN_42121 | _GEN_30332; // @[rob.scala 170:{52,52}]
  wire  _GEN_32575 = _GEN_42122 | _GEN_30333; // @[rob.scala 170:{52,52}]
  wire  _GEN_32576 = _GEN_42123 | _GEN_30334; // @[rob.scala 170:{52,52}]
  wire  _GEN_32577 = _GEN_42124 | _GEN_30335; // @[rob.scala 170:{52,52}]
  wire  _GEN_32578 = _GEN_42125 | _GEN_30336; // @[rob.scala 170:{52,52}]
  wire  _GEN_32579 = _GEN_42126 | _GEN_30337; // @[rob.scala 170:{52,52}]
  wire  _GEN_32580 = _GEN_42127 | _GEN_30338; // @[rob.scala 170:{52,52}]
  wire  _GEN_32581 = _GEN_42128 | _GEN_30339; // @[rob.scala 170:{52,52}]
  wire  _GEN_32582 = io_i_ex_res_packs_0_valid ? _GEN_30406 : _GEN_30212; // @[rob.scala 166:39]
  wire  _GEN_32583 = io_i_ex_res_packs_0_valid ? _GEN_30407 : _GEN_30213; // @[rob.scala 166:39]
  wire  _GEN_32584 = io_i_ex_res_packs_0_valid ? _GEN_30408 : _GEN_30214; // @[rob.scala 166:39]
  wire  _GEN_32585 = io_i_ex_res_packs_0_valid ? _GEN_30409 : _GEN_30215; // @[rob.scala 166:39]
  wire  _GEN_32586 = io_i_ex_res_packs_0_valid ? _GEN_30410 : _GEN_30216; // @[rob.scala 166:39]
  wire  _GEN_32587 = io_i_ex_res_packs_0_valid ? _GEN_30411 : _GEN_30217; // @[rob.scala 166:39]
  wire  _GEN_32588 = io_i_ex_res_packs_0_valid ? _GEN_30412 : _GEN_30218; // @[rob.scala 166:39]
  wire  _GEN_32589 = io_i_ex_res_packs_0_valid ? _GEN_30413 : _GEN_30219; // @[rob.scala 166:39]
  wire  _GEN_32590 = io_i_ex_res_packs_0_valid ? _GEN_30414 : _GEN_30220; // @[rob.scala 166:39]
  wire  _GEN_32591 = io_i_ex_res_packs_0_valid ? _GEN_30415 : _GEN_30221; // @[rob.scala 166:39]
  wire  _GEN_32592 = io_i_ex_res_packs_0_valid ? _GEN_30416 : _GEN_30222; // @[rob.scala 166:39]
  wire  _GEN_32593 = io_i_ex_res_packs_0_valid ? _GEN_30417 : _GEN_30223; // @[rob.scala 166:39]
  wire  _GEN_32594 = io_i_ex_res_packs_0_valid ? _GEN_30418 : _GEN_30224; // @[rob.scala 166:39]
  wire  _GEN_32595 = io_i_ex_res_packs_0_valid ? _GEN_30419 : _GEN_30225; // @[rob.scala 166:39]
  wire  _GEN_32596 = io_i_ex_res_packs_0_valid ? _GEN_30420 : _GEN_30226; // @[rob.scala 166:39]
  wire  _GEN_32597 = io_i_ex_res_packs_0_valid ? _GEN_30421 : _GEN_30227; // @[rob.scala 166:39]
  wire  _GEN_32598 = io_i_ex_res_packs_0_valid ? _GEN_30422 : _GEN_30228; // @[rob.scala 166:39]
  wire  _GEN_32599 = io_i_ex_res_packs_0_valid ? _GEN_30423 : _GEN_30229; // @[rob.scala 166:39]
  wire  _GEN_32600 = io_i_ex_res_packs_0_valid ? _GEN_30424 : _GEN_30230; // @[rob.scala 166:39]
  wire  _GEN_32601 = io_i_ex_res_packs_0_valid ? _GEN_30425 : _GEN_30231; // @[rob.scala 166:39]
  wire  _GEN_32602 = io_i_ex_res_packs_0_valid ? _GEN_30426 : _GEN_30232; // @[rob.scala 166:39]
  wire  _GEN_32603 = io_i_ex_res_packs_0_valid ? _GEN_30427 : _GEN_30233; // @[rob.scala 166:39]
  wire  _GEN_32604 = io_i_ex_res_packs_0_valid ? _GEN_30428 : _GEN_30234; // @[rob.scala 166:39]
  wire  _GEN_32605 = io_i_ex_res_packs_0_valid ? _GEN_30429 : _GEN_30235; // @[rob.scala 166:39]
  wire  _GEN_32606 = io_i_ex_res_packs_0_valid ? _GEN_30430 : _GEN_30236; // @[rob.scala 166:39]
  wire  _GEN_32607 = io_i_ex_res_packs_0_valid ? _GEN_30431 : _GEN_30237; // @[rob.scala 166:39]
  wire  _GEN_32608 = io_i_ex_res_packs_0_valid ? _GEN_30432 : _GEN_30238; // @[rob.scala 166:39]
  wire  _GEN_32609 = io_i_ex_res_packs_0_valid ? _GEN_30433 : _GEN_30239; // @[rob.scala 166:39]
  wire  _GEN_32610 = io_i_ex_res_packs_0_valid ? _GEN_30434 : _GEN_30240; // @[rob.scala 166:39]
  wire  _GEN_32611 = io_i_ex_res_packs_0_valid ? _GEN_30435 : _GEN_30241; // @[rob.scala 166:39]
  wire  _GEN_32612 = io_i_ex_res_packs_0_valid ? _GEN_30436 : _GEN_30242; // @[rob.scala 166:39]
  wire  _GEN_32613 = io_i_ex_res_packs_0_valid ? _GEN_30437 : _GEN_30243; // @[rob.scala 166:39]
  wire  _GEN_32614 = io_i_ex_res_packs_0_valid ? _GEN_30438 : _GEN_30244; // @[rob.scala 166:39]
  wire  _GEN_32615 = io_i_ex_res_packs_0_valid ? _GEN_30439 : _GEN_30245; // @[rob.scala 166:39]
  wire  _GEN_32616 = io_i_ex_res_packs_0_valid ? _GEN_30440 : _GEN_30246; // @[rob.scala 166:39]
  wire  _GEN_32617 = io_i_ex_res_packs_0_valid ? _GEN_30441 : _GEN_30247; // @[rob.scala 166:39]
  wire  _GEN_32618 = io_i_ex_res_packs_0_valid ? _GEN_30442 : _GEN_30248; // @[rob.scala 166:39]
  wire  _GEN_32619 = io_i_ex_res_packs_0_valid ? _GEN_30443 : _GEN_30249; // @[rob.scala 166:39]
  wire  _GEN_32620 = io_i_ex_res_packs_0_valid ? _GEN_30444 : _GEN_30250; // @[rob.scala 166:39]
  wire  _GEN_32621 = io_i_ex_res_packs_0_valid ? _GEN_30445 : _GEN_30251; // @[rob.scala 166:39]
  wire  _GEN_32622 = io_i_ex_res_packs_0_valid ? _GEN_30446 : _GEN_30252; // @[rob.scala 166:39]
  wire  _GEN_32623 = io_i_ex_res_packs_0_valid ? _GEN_30447 : _GEN_30253; // @[rob.scala 166:39]
  wire  _GEN_32624 = io_i_ex_res_packs_0_valid ? _GEN_30448 : _GEN_30254; // @[rob.scala 166:39]
  wire  _GEN_32625 = io_i_ex_res_packs_0_valid ? _GEN_30449 : _GEN_30255; // @[rob.scala 166:39]
  wire  _GEN_32626 = io_i_ex_res_packs_0_valid ? _GEN_30450 : _GEN_30256; // @[rob.scala 166:39]
  wire  _GEN_32627 = io_i_ex_res_packs_0_valid ? _GEN_30451 : _GEN_30257; // @[rob.scala 166:39]
  wire  _GEN_32628 = io_i_ex_res_packs_0_valid ? _GEN_30452 : _GEN_30258; // @[rob.scala 166:39]
  wire  _GEN_32629 = io_i_ex_res_packs_0_valid ? _GEN_30453 : _GEN_30259; // @[rob.scala 166:39]
  wire  _GEN_32630 = io_i_ex_res_packs_0_valid ? _GEN_30454 : _GEN_30260; // @[rob.scala 166:39]
  wire  _GEN_32631 = io_i_ex_res_packs_0_valid ? _GEN_30455 : _GEN_30261; // @[rob.scala 166:39]
  wire  _GEN_32632 = io_i_ex_res_packs_0_valid ? _GEN_30456 : _GEN_30262; // @[rob.scala 166:39]
  wire  _GEN_32633 = io_i_ex_res_packs_0_valid ? _GEN_30457 : _GEN_30263; // @[rob.scala 166:39]
  wire  _GEN_32634 = io_i_ex_res_packs_0_valid ? _GEN_30458 : _GEN_30264; // @[rob.scala 166:39]
  wire  _GEN_32635 = io_i_ex_res_packs_0_valid ? _GEN_30459 : _GEN_30265; // @[rob.scala 166:39]
  wire  _GEN_32636 = io_i_ex_res_packs_0_valid ? _GEN_30460 : _GEN_30266; // @[rob.scala 166:39]
  wire  _GEN_32637 = io_i_ex_res_packs_0_valid ? _GEN_30461 : _GEN_30267; // @[rob.scala 166:39]
  wire  _GEN_32638 = io_i_ex_res_packs_0_valid ? _GEN_30462 : _GEN_30268; // @[rob.scala 166:39]
  wire  _GEN_32639 = io_i_ex_res_packs_0_valid ? _GEN_30463 : _GEN_30269; // @[rob.scala 166:39]
  wire  _GEN_32640 = io_i_ex_res_packs_0_valid ? _GEN_30464 : _GEN_30270; // @[rob.scala 166:39]
  wire  _GEN_32641 = io_i_ex_res_packs_0_valid ? _GEN_30465 : _GEN_30271; // @[rob.scala 166:39]
  wire  _GEN_32642 = io_i_ex_res_packs_0_valid ? _GEN_30466 : _GEN_30272; // @[rob.scala 166:39]
  wire  _GEN_32643 = io_i_ex_res_packs_0_valid ? _GEN_30467 : _GEN_30273; // @[rob.scala 166:39]
  wire  _GEN_32644 = io_i_ex_res_packs_0_valid ? _GEN_30468 : _GEN_30274; // @[rob.scala 166:39]
  wire  _GEN_32645 = io_i_ex_res_packs_0_valid ? _GEN_30469 : _GEN_30275; // @[rob.scala 166:39]
  wire [31:0] _GEN_32710 = io_i_ex_res_packs_0_valid ? _GEN_30534 : _GEN_28292; // @[rob.scala 166:39]
  wire [31:0] _GEN_32711 = io_i_ex_res_packs_0_valid ? _GEN_30535 : _GEN_28293; // @[rob.scala 166:39]
  wire [31:0] _GEN_32712 = io_i_ex_res_packs_0_valid ? _GEN_30536 : _GEN_28294; // @[rob.scala 166:39]
  wire [31:0] _GEN_32713 = io_i_ex_res_packs_0_valid ? _GEN_30537 : _GEN_28295; // @[rob.scala 166:39]
  wire [31:0] _GEN_32714 = io_i_ex_res_packs_0_valid ? _GEN_30538 : _GEN_28296; // @[rob.scala 166:39]
  wire [31:0] _GEN_32715 = io_i_ex_res_packs_0_valid ? _GEN_30539 : _GEN_28297; // @[rob.scala 166:39]
  wire [31:0] _GEN_32716 = io_i_ex_res_packs_0_valid ? _GEN_30540 : _GEN_28298; // @[rob.scala 166:39]
  wire [31:0] _GEN_32717 = io_i_ex_res_packs_0_valid ? _GEN_30541 : _GEN_28299; // @[rob.scala 166:39]
  wire [31:0] _GEN_32718 = io_i_ex_res_packs_0_valid ? _GEN_30542 : _GEN_28300; // @[rob.scala 166:39]
  wire [31:0] _GEN_32719 = io_i_ex_res_packs_0_valid ? _GEN_30543 : _GEN_28301; // @[rob.scala 166:39]
  wire [31:0] _GEN_32720 = io_i_ex_res_packs_0_valid ? _GEN_30544 : _GEN_28302; // @[rob.scala 166:39]
  wire [31:0] _GEN_32721 = io_i_ex_res_packs_0_valid ? _GEN_30545 : _GEN_28303; // @[rob.scala 166:39]
  wire [31:0] _GEN_32722 = io_i_ex_res_packs_0_valid ? _GEN_30546 : _GEN_28304; // @[rob.scala 166:39]
  wire [31:0] _GEN_32723 = io_i_ex_res_packs_0_valid ? _GEN_30547 : _GEN_28305; // @[rob.scala 166:39]
  wire [31:0] _GEN_32724 = io_i_ex_res_packs_0_valid ? _GEN_30548 : _GEN_28306; // @[rob.scala 166:39]
  wire [31:0] _GEN_32725 = io_i_ex_res_packs_0_valid ? _GEN_30549 : _GEN_28307; // @[rob.scala 166:39]
  wire [31:0] _GEN_32726 = io_i_ex_res_packs_0_valid ? _GEN_30550 : _GEN_28308; // @[rob.scala 166:39]
  wire [31:0] _GEN_32727 = io_i_ex_res_packs_0_valid ? _GEN_30551 : _GEN_28309; // @[rob.scala 166:39]
  wire [31:0] _GEN_32728 = io_i_ex_res_packs_0_valid ? _GEN_30552 : _GEN_28310; // @[rob.scala 166:39]
  wire [31:0] _GEN_32729 = io_i_ex_res_packs_0_valid ? _GEN_30553 : _GEN_28311; // @[rob.scala 166:39]
  wire [31:0] _GEN_32730 = io_i_ex_res_packs_0_valid ? _GEN_30554 : _GEN_28312; // @[rob.scala 166:39]
  wire [31:0] _GEN_32731 = io_i_ex_res_packs_0_valid ? _GEN_30555 : _GEN_28313; // @[rob.scala 166:39]
  wire [31:0] _GEN_32732 = io_i_ex_res_packs_0_valid ? _GEN_30556 : _GEN_28314; // @[rob.scala 166:39]
  wire [31:0] _GEN_32733 = io_i_ex_res_packs_0_valid ? _GEN_30557 : _GEN_28315; // @[rob.scala 166:39]
  wire [31:0] _GEN_32734 = io_i_ex_res_packs_0_valid ? _GEN_30558 : _GEN_28316; // @[rob.scala 166:39]
  wire [31:0] _GEN_32735 = io_i_ex_res_packs_0_valid ? _GEN_30559 : _GEN_28317; // @[rob.scala 166:39]
  wire [31:0] _GEN_32736 = io_i_ex_res_packs_0_valid ? _GEN_30560 : _GEN_28318; // @[rob.scala 166:39]
  wire [31:0] _GEN_32737 = io_i_ex_res_packs_0_valid ? _GEN_30561 : _GEN_28319; // @[rob.scala 166:39]
  wire [31:0] _GEN_32738 = io_i_ex_res_packs_0_valid ? _GEN_30562 : _GEN_28320; // @[rob.scala 166:39]
  wire [31:0] _GEN_32739 = io_i_ex_res_packs_0_valid ? _GEN_30563 : _GEN_28321; // @[rob.scala 166:39]
  wire [31:0] _GEN_32740 = io_i_ex_res_packs_0_valid ? _GEN_30564 : _GEN_28322; // @[rob.scala 166:39]
  wire [31:0] _GEN_32741 = io_i_ex_res_packs_0_valid ? _GEN_30565 : _GEN_28323; // @[rob.scala 166:39]
  wire [31:0] _GEN_32742 = io_i_ex_res_packs_0_valid ? _GEN_30566 : _GEN_28324; // @[rob.scala 166:39]
  wire [31:0] _GEN_32743 = io_i_ex_res_packs_0_valid ? _GEN_30567 : _GEN_28325; // @[rob.scala 166:39]
  wire [31:0] _GEN_32744 = io_i_ex_res_packs_0_valid ? _GEN_30568 : _GEN_28326; // @[rob.scala 166:39]
  wire [31:0] _GEN_32745 = io_i_ex_res_packs_0_valid ? _GEN_30569 : _GEN_28327; // @[rob.scala 166:39]
  wire [31:0] _GEN_32746 = io_i_ex_res_packs_0_valid ? _GEN_30570 : _GEN_28328; // @[rob.scala 166:39]
  wire [31:0] _GEN_32747 = io_i_ex_res_packs_0_valid ? _GEN_30571 : _GEN_28329; // @[rob.scala 166:39]
  wire [31:0] _GEN_32748 = io_i_ex_res_packs_0_valid ? _GEN_30572 : _GEN_28330; // @[rob.scala 166:39]
  wire [31:0] _GEN_32749 = io_i_ex_res_packs_0_valid ? _GEN_30573 : _GEN_28331; // @[rob.scala 166:39]
  wire [31:0] _GEN_32750 = io_i_ex_res_packs_0_valid ? _GEN_30574 : _GEN_28332; // @[rob.scala 166:39]
  wire [31:0] _GEN_32751 = io_i_ex_res_packs_0_valid ? _GEN_30575 : _GEN_28333; // @[rob.scala 166:39]
  wire [31:0] _GEN_32752 = io_i_ex_res_packs_0_valid ? _GEN_30576 : _GEN_28334; // @[rob.scala 166:39]
  wire [31:0] _GEN_32753 = io_i_ex_res_packs_0_valid ? _GEN_30577 : _GEN_28335; // @[rob.scala 166:39]
  wire [31:0] _GEN_32754 = io_i_ex_res_packs_0_valid ? _GEN_30578 : _GEN_28336; // @[rob.scala 166:39]
  wire [31:0] _GEN_32755 = io_i_ex_res_packs_0_valid ? _GEN_30579 : _GEN_28337; // @[rob.scala 166:39]
  wire [31:0] _GEN_32756 = io_i_ex_res_packs_0_valid ? _GEN_30580 : _GEN_28338; // @[rob.scala 166:39]
  wire [31:0] _GEN_32757 = io_i_ex_res_packs_0_valid ? _GEN_30581 : _GEN_28339; // @[rob.scala 166:39]
  wire [31:0] _GEN_32758 = io_i_ex_res_packs_0_valid ? _GEN_30582 : _GEN_28340; // @[rob.scala 166:39]
  wire [31:0] _GEN_32759 = io_i_ex_res_packs_0_valid ? _GEN_30583 : _GEN_28341; // @[rob.scala 166:39]
  wire [31:0] _GEN_32760 = io_i_ex_res_packs_0_valid ? _GEN_30584 : _GEN_28342; // @[rob.scala 166:39]
  wire [31:0] _GEN_32761 = io_i_ex_res_packs_0_valid ? _GEN_30585 : _GEN_28343; // @[rob.scala 166:39]
  wire [31:0] _GEN_32762 = io_i_ex_res_packs_0_valid ? _GEN_30586 : _GEN_28344; // @[rob.scala 166:39]
  wire [31:0] _GEN_32763 = io_i_ex_res_packs_0_valid ? _GEN_30587 : _GEN_28345; // @[rob.scala 166:39]
  wire [31:0] _GEN_32764 = io_i_ex_res_packs_0_valid ? _GEN_30588 : _GEN_28346; // @[rob.scala 166:39]
  wire [31:0] _GEN_32765 = io_i_ex_res_packs_0_valid ? _GEN_30589 : _GEN_28347; // @[rob.scala 166:39]
  wire [31:0] _GEN_32766 = io_i_ex_res_packs_0_valid ? _GEN_30590 : _GEN_28348; // @[rob.scala 166:39]
  wire [31:0] _GEN_32767 = io_i_ex_res_packs_0_valid ? _GEN_30591 : _GEN_28349; // @[rob.scala 166:39]
  wire [31:0] _GEN_32768 = io_i_ex_res_packs_0_valid ? _GEN_30592 : _GEN_28350; // @[rob.scala 166:39]
  wire [31:0] _GEN_32769 = io_i_ex_res_packs_0_valid ? _GEN_30593 : _GEN_28351; // @[rob.scala 166:39]
  wire [31:0] _GEN_32770 = io_i_ex_res_packs_0_valid ? _GEN_30594 : _GEN_28352; // @[rob.scala 166:39]
  wire [31:0] _GEN_32771 = io_i_ex_res_packs_0_valid ? _GEN_30595 : _GEN_28353; // @[rob.scala 166:39]
  wire [31:0] _GEN_32772 = io_i_ex_res_packs_0_valid ? _GEN_30596 : _GEN_28354; // @[rob.scala 166:39]
  wire [31:0] _GEN_32773 = io_i_ex_res_packs_0_valid ? _GEN_30597 : _GEN_28355; // @[rob.scala 166:39]
  wire [31:0] _GEN_32774 = io_i_ex_res_packs_0_valid ? _GEN_30598 : _GEN_28356; // @[rob.scala 166:39]
  wire [31:0] _GEN_32775 = io_i_ex_res_packs_0_valid ? _GEN_30599 : _GEN_28357; // @[rob.scala 166:39]
  wire [31:0] _GEN_32776 = io_i_ex_res_packs_0_valid ? _GEN_30600 : _GEN_28358; // @[rob.scala 166:39]
  wire [31:0] _GEN_32777 = io_i_ex_res_packs_0_valid ? _GEN_30601 : _GEN_28359; // @[rob.scala 166:39]
  wire [31:0] _GEN_32778 = io_i_ex_res_packs_0_valid ? _GEN_30602 : _GEN_28360; // @[rob.scala 166:39]
  wire [31:0] _GEN_32779 = io_i_ex_res_packs_0_valid ? _GEN_30603 : _GEN_28361; // @[rob.scala 166:39]
  wire [31:0] _GEN_32780 = io_i_ex_res_packs_0_valid ? _GEN_30604 : _GEN_28362; // @[rob.scala 166:39]
  wire [31:0] _GEN_32781 = io_i_ex_res_packs_0_valid ? _GEN_30605 : _GEN_28363; // @[rob.scala 166:39]
  wire [31:0] _GEN_32782 = io_i_ex_res_packs_0_valid ? _GEN_30606 : _GEN_28364; // @[rob.scala 166:39]
  wire [31:0] _GEN_32783 = io_i_ex_res_packs_0_valid ? _GEN_30607 : _GEN_28365; // @[rob.scala 166:39]
  wire [31:0] _GEN_32784 = io_i_ex_res_packs_0_valid ? _GEN_30608 : _GEN_28366; // @[rob.scala 166:39]
  wire [31:0] _GEN_32785 = io_i_ex_res_packs_0_valid ? _GEN_30609 : _GEN_28367; // @[rob.scala 166:39]
  wire [31:0] _GEN_32786 = io_i_ex_res_packs_0_valid ? _GEN_30610 : _GEN_28368; // @[rob.scala 166:39]
  wire [31:0] _GEN_32787 = io_i_ex_res_packs_0_valid ? _GEN_30611 : _GEN_28369; // @[rob.scala 166:39]
  wire [31:0] _GEN_32788 = io_i_ex_res_packs_0_valid ? _GEN_30612 : _GEN_28370; // @[rob.scala 166:39]
  wire [31:0] _GEN_32789 = io_i_ex_res_packs_0_valid ? _GEN_30613 : _GEN_28371; // @[rob.scala 166:39]
  wire [31:0] _GEN_32790 = io_i_ex_res_packs_0_valid ? _GEN_30614 : _GEN_28372; // @[rob.scala 166:39]
  wire [31:0] _GEN_32791 = io_i_ex_res_packs_0_valid ? _GEN_30615 : _GEN_28373; // @[rob.scala 166:39]
  wire [31:0] _GEN_32792 = io_i_ex_res_packs_0_valid ? _GEN_30616 : _GEN_28374; // @[rob.scala 166:39]
  wire [31:0] _GEN_32793 = io_i_ex_res_packs_0_valid ? _GEN_30617 : _GEN_28375; // @[rob.scala 166:39]
  wire [31:0] _GEN_32794 = io_i_ex_res_packs_0_valid ? _GEN_30618 : _GEN_28376; // @[rob.scala 166:39]
  wire [31:0] _GEN_32795 = io_i_ex_res_packs_0_valid ? _GEN_30619 : _GEN_28377; // @[rob.scala 166:39]
  wire [31:0] _GEN_32796 = io_i_ex_res_packs_0_valid ? _GEN_30620 : _GEN_28378; // @[rob.scala 166:39]
  wire [31:0] _GEN_32797 = io_i_ex_res_packs_0_valid ? _GEN_30621 : _GEN_28379; // @[rob.scala 166:39]
  wire [31:0] _GEN_32798 = io_i_ex_res_packs_0_valid ? _GEN_30622 : _GEN_28380; // @[rob.scala 166:39]
  wire [31:0] _GEN_32799 = io_i_ex_res_packs_0_valid ? _GEN_30623 : _GEN_28381; // @[rob.scala 166:39]
  wire [31:0] _GEN_32800 = io_i_ex_res_packs_0_valid ? _GEN_30624 : _GEN_28382; // @[rob.scala 166:39]
  wire [31:0] _GEN_32801 = io_i_ex_res_packs_0_valid ? _GEN_30625 : _GEN_28383; // @[rob.scala 166:39]
  wire [31:0] _GEN_32802 = io_i_ex_res_packs_0_valid ? _GEN_30626 : _GEN_28384; // @[rob.scala 166:39]
  wire [31:0] _GEN_32803 = io_i_ex_res_packs_0_valid ? _GEN_30627 : _GEN_28385; // @[rob.scala 166:39]
  wire [31:0] _GEN_32804 = io_i_ex_res_packs_0_valid ? _GEN_30628 : _GEN_28386; // @[rob.scala 166:39]
  wire [31:0] _GEN_32805 = io_i_ex_res_packs_0_valid ? _GEN_30629 : _GEN_28387; // @[rob.scala 166:39]
  wire [31:0] _GEN_32806 = io_i_ex_res_packs_0_valid ? _GEN_30630 : _GEN_28388; // @[rob.scala 166:39]
  wire [31:0] _GEN_32807 = io_i_ex_res_packs_0_valid ? _GEN_30631 : _GEN_28389; // @[rob.scala 166:39]
  wire [31:0] _GEN_32808 = io_i_ex_res_packs_0_valid ? _GEN_30632 : _GEN_28390; // @[rob.scala 166:39]
  wire [31:0] _GEN_32809 = io_i_ex_res_packs_0_valid ? _GEN_30633 : _GEN_28391; // @[rob.scala 166:39]
  wire [31:0] _GEN_32810 = io_i_ex_res_packs_0_valid ? _GEN_30634 : _GEN_28392; // @[rob.scala 166:39]
  wire [31:0] _GEN_32811 = io_i_ex_res_packs_0_valid ? _GEN_30635 : _GEN_28393; // @[rob.scala 166:39]
  wire [31:0] _GEN_32812 = io_i_ex_res_packs_0_valid ? _GEN_30636 : _GEN_28394; // @[rob.scala 166:39]
  wire [31:0] _GEN_32813 = io_i_ex_res_packs_0_valid ? _GEN_30637 : _GEN_28395; // @[rob.scala 166:39]
  wire [31:0] _GEN_32814 = io_i_ex_res_packs_0_valid ? _GEN_30638 : _GEN_28396; // @[rob.scala 166:39]
  wire [31:0] _GEN_32815 = io_i_ex_res_packs_0_valid ? _GEN_30639 : _GEN_28397; // @[rob.scala 166:39]
  wire [31:0] _GEN_32816 = io_i_ex_res_packs_0_valid ? _GEN_30640 : _GEN_28398; // @[rob.scala 166:39]
  wire [31:0] _GEN_32817 = io_i_ex_res_packs_0_valid ? _GEN_30641 : _GEN_28399; // @[rob.scala 166:39]
  wire [31:0] _GEN_32818 = io_i_ex_res_packs_0_valid ? _GEN_30642 : _GEN_28400; // @[rob.scala 166:39]
  wire [31:0] _GEN_32819 = io_i_ex_res_packs_0_valid ? _GEN_30643 : _GEN_28401; // @[rob.scala 166:39]
  wire [31:0] _GEN_32820 = io_i_ex_res_packs_0_valid ? _GEN_30644 : _GEN_28402; // @[rob.scala 166:39]
  wire [31:0] _GEN_32821 = io_i_ex_res_packs_0_valid ? _GEN_30645 : _GEN_28403; // @[rob.scala 166:39]
  wire [31:0] _GEN_32822 = io_i_ex_res_packs_0_valid ? _GEN_30646 : _GEN_28404; // @[rob.scala 166:39]
  wire [31:0] _GEN_32823 = io_i_ex_res_packs_0_valid ? _GEN_30647 : _GEN_28405; // @[rob.scala 166:39]
  wire [31:0] _GEN_32824 = io_i_ex_res_packs_0_valid ? _GEN_30648 : _GEN_28406; // @[rob.scala 166:39]
  wire [31:0] _GEN_32825 = io_i_ex_res_packs_0_valid ? _GEN_30649 : _GEN_28407; // @[rob.scala 166:39]
  wire [31:0] _GEN_32826 = io_i_ex_res_packs_0_valid ? _GEN_30650 : _GEN_28408; // @[rob.scala 166:39]
  wire [31:0] _GEN_32827 = io_i_ex_res_packs_0_valid ? _GEN_30651 : _GEN_28409; // @[rob.scala 166:39]
  wire [31:0] _GEN_32828 = io_i_ex_res_packs_0_valid ? _GEN_30652 : _GEN_28410; // @[rob.scala 166:39]
  wire [31:0] _GEN_32829 = io_i_ex_res_packs_0_valid ? _GEN_30653 : _GEN_28411; // @[rob.scala 166:39]
  wire [31:0] _GEN_32830 = io_i_ex_res_packs_0_valid ? _GEN_30654 : _GEN_28412; // @[rob.scala 166:39]
  wire [31:0] _GEN_32831 = io_i_ex_res_packs_0_valid ? _GEN_30655 : _GEN_28413; // @[rob.scala 166:39]
  wire [31:0] _GEN_32832 = io_i_ex_res_packs_0_valid ? _GEN_30656 : _GEN_28414; // @[rob.scala 166:39]
  wire [31:0] _GEN_32833 = io_i_ex_res_packs_0_valid ? _GEN_30657 : _GEN_28415; // @[rob.scala 166:39]
  wire [31:0] _GEN_32834 = io_i_ex_res_packs_0_valid ? _GEN_30658 : _GEN_28416; // @[rob.scala 166:39]
  wire [31:0] _GEN_32835 = io_i_ex_res_packs_0_valid ? _GEN_30659 : _GEN_28417; // @[rob.scala 166:39]
  wire [31:0] _GEN_32836 = io_i_ex_res_packs_0_valid ? _GEN_30660 : _GEN_28418; // @[rob.scala 166:39]
  wire [31:0] _GEN_32837 = io_i_ex_res_packs_0_valid ? _GEN_30661 : _GEN_28419; // @[rob.scala 166:39]
  wire [6:0] _GEN_32838 = io_i_ex_res_packs_0_valid ? _GEN_30662 : _GEN_28420; // @[rob.scala 166:39]
  wire [6:0] _GEN_32839 = io_i_ex_res_packs_0_valid ? _GEN_30663 : _GEN_28421; // @[rob.scala 166:39]
  wire [6:0] _GEN_32840 = io_i_ex_res_packs_0_valid ? _GEN_30664 : _GEN_28422; // @[rob.scala 166:39]
  wire [6:0] _GEN_32841 = io_i_ex_res_packs_0_valid ? _GEN_30665 : _GEN_28423; // @[rob.scala 166:39]
  wire [6:0] _GEN_32842 = io_i_ex_res_packs_0_valid ? _GEN_30666 : _GEN_28424; // @[rob.scala 166:39]
  wire [6:0] _GEN_32843 = io_i_ex_res_packs_0_valid ? _GEN_30667 : _GEN_28425; // @[rob.scala 166:39]
  wire [6:0] _GEN_32844 = io_i_ex_res_packs_0_valid ? _GEN_30668 : _GEN_28426; // @[rob.scala 166:39]
  wire [6:0] _GEN_32845 = io_i_ex_res_packs_0_valid ? _GEN_30669 : _GEN_28427; // @[rob.scala 166:39]
  wire [6:0] _GEN_32846 = io_i_ex_res_packs_0_valid ? _GEN_30670 : _GEN_28428; // @[rob.scala 166:39]
  wire [6:0] _GEN_32847 = io_i_ex_res_packs_0_valid ? _GEN_30671 : _GEN_28429; // @[rob.scala 166:39]
  wire [6:0] _GEN_32848 = io_i_ex_res_packs_0_valid ? _GEN_30672 : _GEN_28430; // @[rob.scala 166:39]
  wire [6:0] _GEN_32849 = io_i_ex_res_packs_0_valid ? _GEN_30673 : _GEN_28431; // @[rob.scala 166:39]
  wire [6:0] _GEN_32850 = io_i_ex_res_packs_0_valid ? _GEN_30674 : _GEN_28432; // @[rob.scala 166:39]
  wire [6:0] _GEN_32851 = io_i_ex_res_packs_0_valid ? _GEN_30675 : _GEN_28433; // @[rob.scala 166:39]
  wire [6:0] _GEN_32852 = io_i_ex_res_packs_0_valid ? _GEN_30676 : _GEN_28434; // @[rob.scala 166:39]
  wire [6:0] _GEN_32853 = io_i_ex_res_packs_0_valid ? _GEN_30677 : _GEN_28435; // @[rob.scala 166:39]
  wire [6:0] _GEN_32854 = io_i_ex_res_packs_0_valid ? _GEN_30678 : _GEN_28436; // @[rob.scala 166:39]
  wire [6:0] _GEN_32855 = io_i_ex_res_packs_0_valid ? _GEN_30679 : _GEN_28437; // @[rob.scala 166:39]
  wire [6:0] _GEN_32856 = io_i_ex_res_packs_0_valid ? _GEN_30680 : _GEN_28438; // @[rob.scala 166:39]
  wire [6:0] _GEN_32857 = io_i_ex_res_packs_0_valid ? _GEN_30681 : _GEN_28439; // @[rob.scala 166:39]
  wire [6:0] _GEN_32858 = io_i_ex_res_packs_0_valid ? _GEN_30682 : _GEN_28440; // @[rob.scala 166:39]
  wire [6:0] _GEN_32859 = io_i_ex_res_packs_0_valid ? _GEN_30683 : _GEN_28441; // @[rob.scala 166:39]
  wire [6:0] _GEN_32860 = io_i_ex_res_packs_0_valid ? _GEN_30684 : _GEN_28442; // @[rob.scala 166:39]
  wire [6:0] _GEN_32861 = io_i_ex_res_packs_0_valid ? _GEN_30685 : _GEN_28443; // @[rob.scala 166:39]
  wire [6:0] _GEN_32862 = io_i_ex_res_packs_0_valid ? _GEN_30686 : _GEN_28444; // @[rob.scala 166:39]
  wire [6:0] _GEN_32863 = io_i_ex_res_packs_0_valid ? _GEN_30687 : _GEN_28445; // @[rob.scala 166:39]
  wire [6:0] _GEN_32864 = io_i_ex_res_packs_0_valid ? _GEN_30688 : _GEN_28446; // @[rob.scala 166:39]
  wire [6:0] _GEN_32865 = io_i_ex_res_packs_0_valid ? _GEN_30689 : _GEN_28447; // @[rob.scala 166:39]
  wire [6:0] _GEN_32866 = io_i_ex_res_packs_0_valid ? _GEN_30690 : _GEN_28448; // @[rob.scala 166:39]
  wire [6:0] _GEN_32867 = io_i_ex_res_packs_0_valid ? _GEN_30691 : _GEN_28449; // @[rob.scala 166:39]
  wire [6:0] _GEN_32868 = io_i_ex_res_packs_0_valid ? _GEN_30692 : _GEN_28450; // @[rob.scala 166:39]
  wire [6:0] _GEN_32869 = io_i_ex_res_packs_0_valid ? _GEN_30693 : _GEN_28451; // @[rob.scala 166:39]
  wire [6:0] _GEN_32870 = io_i_ex_res_packs_0_valid ? _GEN_30694 : _GEN_28452; // @[rob.scala 166:39]
  wire [6:0] _GEN_32871 = io_i_ex_res_packs_0_valid ? _GEN_30695 : _GEN_28453; // @[rob.scala 166:39]
  wire [6:0] _GEN_32872 = io_i_ex_res_packs_0_valid ? _GEN_30696 : _GEN_28454; // @[rob.scala 166:39]
  wire [6:0] _GEN_32873 = io_i_ex_res_packs_0_valid ? _GEN_30697 : _GEN_28455; // @[rob.scala 166:39]
  wire [6:0] _GEN_32874 = io_i_ex_res_packs_0_valid ? _GEN_30698 : _GEN_28456; // @[rob.scala 166:39]
  wire [6:0] _GEN_32875 = io_i_ex_res_packs_0_valid ? _GEN_30699 : _GEN_28457; // @[rob.scala 166:39]
  wire [6:0] _GEN_32876 = io_i_ex_res_packs_0_valid ? _GEN_30700 : _GEN_28458; // @[rob.scala 166:39]
  wire [6:0] _GEN_32877 = io_i_ex_res_packs_0_valid ? _GEN_30701 : _GEN_28459; // @[rob.scala 166:39]
  wire [6:0] _GEN_32878 = io_i_ex_res_packs_0_valid ? _GEN_30702 : _GEN_28460; // @[rob.scala 166:39]
  wire [6:0] _GEN_32879 = io_i_ex_res_packs_0_valid ? _GEN_30703 : _GEN_28461; // @[rob.scala 166:39]
  wire [6:0] _GEN_32880 = io_i_ex_res_packs_0_valid ? _GEN_30704 : _GEN_28462; // @[rob.scala 166:39]
  wire [6:0] _GEN_32881 = io_i_ex_res_packs_0_valid ? _GEN_30705 : _GEN_28463; // @[rob.scala 166:39]
  wire [6:0] _GEN_32882 = io_i_ex_res_packs_0_valid ? _GEN_30706 : _GEN_28464; // @[rob.scala 166:39]
  wire [6:0] _GEN_32883 = io_i_ex_res_packs_0_valid ? _GEN_30707 : _GEN_28465; // @[rob.scala 166:39]
  wire [6:0] _GEN_32884 = io_i_ex_res_packs_0_valid ? _GEN_30708 : _GEN_28466; // @[rob.scala 166:39]
  wire [6:0] _GEN_32885 = io_i_ex_res_packs_0_valid ? _GEN_30709 : _GEN_28467; // @[rob.scala 166:39]
  wire [6:0] _GEN_32886 = io_i_ex_res_packs_0_valid ? _GEN_30710 : _GEN_28468; // @[rob.scala 166:39]
  wire [6:0] _GEN_32887 = io_i_ex_res_packs_0_valid ? _GEN_30711 : _GEN_28469; // @[rob.scala 166:39]
  wire [6:0] _GEN_32888 = io_i_ex_res_packs_0_valid ? _GEN_30712 : _GEN_28470; // @[rob.scala 166:39]
  wire [6:0] _GEN_32889 = io_i_ex_res_packs_0_valid ? _GEN_30713 : _GEN_28471; // @[rob.scala 166:39]
  wire [6:0] _GEN_32890 = io_i_ex_res_packs_0_valid ? _GEN_30714 : _GEN_28472; // @[rob.scala 166:39]
  wire [6:0] _GEN_32891 = io_i_ex_res_packs_0_valid ? _GEN_30715 : _GEN_28473; // @[rob.scala 166:39]
  wire [6:0] _GEN_32892 = io_i_ex_res_packs_0_valid ? _GEN_30716 : _GEN_28474; // @[rob.scala 166:39]
  wire [6:0] _GEN_32893 = io_i_ex_res_packs_0_valid ? _GEN_30717 : _GEN_28475; // @[rob.scala 166:39]
  wire [6:0] _GEN_32894 = io_i_ex_res_packs_0_valid ? _GEN_30718 : _GEN_28476; // @[rob.scala 166:39]
  wire [6:0] _GEN_32895 = io_i_ex_res_packs_0_valid ? _GEN_30719 : _GEN_28477; // @[rob.scala 166:39]
  wire [6:0] _GEN_32896 = io_i_ex_res_packs_0_valid ? _GEN_30720 : _GEN_28478; // @[rob.scala 166:39]
  wire [6:0] _GEN_32897 = io_i_ex_res_packs_0_valid ? _GEN_30721 : _GEN_28479; // @[rob.scala 166:39]
  wire [6:0] _GEN_32898 = io_i_ex_res_packs_0_valid ? _GEN_30722 : _GEN_28480; // @[rob.scala 166:39]
  wire [6:0] _GEN_32899 = io_i_ex_res_packs_0_valid ? _GEN_30723 : _GEN_28481; // @[rob.scala 166:39]
  wire [6:0] _GEN_32900 = io_i_ex_res_packs_0_valid ? _GEN_30724 : _GEN_28482; // @[rob.scala 166:39]
  wire [6:0] _GEN_32901 = io_i_ex_res_packs_0_valid ? _GEN_30725 : _GEN_28483; // @[rob.scala 166:39]
  wire [6:0] _GEN_33222 = io_i_ex_res_packs_0_valid ? _GEN_31046 : _GEN_28804; // @[rob.scala 166:39]
  wire [6:0] _GEN_33223 = io_i_ex_res_packs_0_valid ? _GEN_31047 : _GEN_28805; // @[rob.scala 166:39]
  wire [6:0] _GEN_33224 = io_i_ex_res_packs_0_valid ? _GEN_31048 : _GEN_28806; // @[rob.scala 166:39]
  wire [6:0] _GEN_33225 = io_i_ex_res_packs_0_valid ? _GEN_31049 : _GEN_28807; // @[rob.scala 166:39]
  wire [6:0] _GEN_33226 = io_i_ex_res_packs_0_valid ? _GEN_31050 : _GEN_28808; // @[rob.scala 166:39]
  wire [6:0] _GEN_33227 = io_i_ex_res_packs_0_valid ? _GEN_31051 : _GEN_28809; // @[rob.scala 166:39]
  wire [6:0] _GEN_33228 = io_i_ex_res_packs_0_valid ? _GEN_31052 : _GEN_28810; // @[rob.scala 166:39]
  wire [6:0] _GEN_33229 = io_i_ex_res_packs_0_valid ? _GEN_31053 : _GEN_28811; // @[rob.scala 166:39]
  wire [6:0] _GEN_33230 = io_i_ex_res_packs_0_valid ? _GEN_31054 : _GEN_28812; // @[rob.scala 166:39]
  wire [6:0] _GEN_33231 = io_i_ex_res_packs_0_valid ? _GEN_31055 : _GEN_28813; // @[rob.scala 166:39]
  wire [6:0] _GEN_33232 = io_i_ex_res_packs_0_valid ? _GEN_31056 : _GEN_28814; // @[rob.scala 166:39]
  wire [6:0] _GEN_33233 = io_i_ex_res_packs_0_valid ? _GEN_31057 : _GEN_28815; // @[rob.scala 166:39]
  wire [6:0] _GEN_33234 = io_i_ex_res_packs_0_valid ? _GEN_31058 : _GEN_28816; // @[rob.scala 166:39]
  wire [6:0] _GEN_33235 = io_i_ex_res_packs_0_valid ? _GEN_31059 : _GEN_28817; // @[rob.scala 166:39]
  wire [6:0] _GEN_33236 = io_i_ex_res_packs_0_valid ? _GEN_31060 : _GEN_28818; // @[rob.scala 166:39]
  wire [6:0] _GEN_33237 = io_i_ex_res_packs_0_valid ? _GEN_31061 : _GEN_28819; // @[rob.scala 166:39]
  wire [6:0] _GEN_33238 = io_i_ex_res_packs_0_valid ? _GEN_31062 : _GEN_28820; // @[rob.scala 166:39]
  wire [6:0] _GEN_33239 = io_i_ex_res_packs_0_valid ? _GEN_31063 : _GEN_28821; // @[rob.scala 166:39]
  wire [6:0] _GEN_33240 = io_i_ex_res_packs_0_valid ? _GEN_31064 : _GEN_28822; // @[rob.scala 166:39]
  wire [6:0] _GEN_33241 = io_i_ex_res_packs_0_valid ? _GEN_31065 : _GEN_28823; // @[rob.scala 166:39]
  wire [6:0] _GEN_33242 = io_i_ex_res_packs_0_valid ? _GEN_31066 : _GEN_28824; // @[rob.scala 166:39]
  wire [6:0] _GEN_33243 = io_i_ex_res_packs_0_valid ? _GEN_31067 : _GEN_28825; // @[rob.scala 166:39]
  wire [6:0] _GEN_33244 = io_i_ex_res_packs_0_valid ? _GEN_31068 : _GEN_28826; // @[rob.scala 166:39]
  wire [6:0] _GEN_33245 = io_i_ex_res_packs_0_valid ? _GEN_31069 : _GEN_28827; // @[rob.scala 166:39]
  wire [6:0] _GEN_33246 = io_i_ex_res_packs_0_valid ? _GEN_31070 : _GEN_28828; // @[rob.scala 166:39]
  wire [6:0] _GEN_33247 = io_i_ex_res_packs_0_valid ? _GEN_31071 : _GEN_28829; // @[rob.scala 166:39]
  wire [6:0] _GEN_33248 = io_i_ex_res_packs_0_valid ? _GEN_31072 : _GEN_28830; // @[rob.scala 166:39]
  wire [6:0] _GEN_33249 = io_i_ex_res_packs_0_valid ? _GEN_31073 : _GEN_28831; // @[rob.scala 166:39]
  wire [6:0] _GEN_33250 = io_i_ex_res_packs_0_valid ? _GEN_31074 : _GEN_28832; // @[rob.scala 166:39]
  wire [6:0] _GEN_33251 = io_i_ex_res_packs_0_valid ? _GEN_31075 : _GEN_28833; // @[rob.scala 166:39]
  wire [6:0] _GEN_33252 = io_i_ex_res_packs_0_valid ? _GEN_31076 : _GEN_28834; // @[rob.scala 166:39]
  wire [6:0] _GEN_33253 = io_i_ex_res_packs_0_valid ? _GEN_31077 : _GEN_28835; // @[rob.scala 166:39]
  wire [6:0] _GEN_33254 = io_i_ex_res_packs_0_valid ? _GEN_31078 : _GEN_28836; // @[rob.scala 166:39]
  wire [6:0] _GEN_33255 = io_i_ex_res_packs_0_valid ? _GEN_31079 : _GEN_28837; // @[rob.scala 166:39]
  wire [6:0] _GEN_33256 = io_i_ex_res_packs_0_valid ? _GEN_31080 : _GEN_28838; // @[rob.scala 166:39]
  wire [6:0] _GEN_33257 = io_i_ex_res_packs_0_valid ? _GEN_31081 : _GEN_28839; // @[rob.scala 166:39]
  wire [6:0] _GEN_33258 = io_i_ex_res_packs_0_valid ? _GEN_31082 : _GEN_28840; // @[rob.scala 166:39]
  wire [6:0] _GEN_33259 = io_i_ex_res_packs_0_valid ? _GEN_31083 : _GEN_28841; // @[rob.scala 166:39]
  wire [6:0] _GEN_33260 = io_i_ex_res_packs_0_valid ? _GEN_31084 : _GEN_28842; // @[rob.scala 166:39]
  wire [6:0] _GEN_33261 = io_i_ex_res_packs_0_valid ? _GEN_31085 : _GEN_28843; // @[rob.scala 166:39]
  wire [6:0] _GEN_33262 = io_i_ex_res_packs_0_valid ? _GEN_31086 : _GEN_28844; // @[rob.scala 166:39]
  wire [6:0] _GEN_33263 = io_i_ex_res_packs_0_valid ? _GEN_31087 : _GEN_28845; // @[rob.scala 166:39]
  wire [6:0] _GEN_33264 = io_i_ex_res_packs_0_valid ? _GEN_31088 : _GEN_28846; // @[rob.scala 166:39]
  wire [6:0] _GEN_33265 = io_i_ex_res_packs_0_valid ? _GEN_31089 : _GEN_28847; // @[rob.scala 166:39]
  wire [6:0] _GEN_33266 = io_i_ex_res_packs_0_valid ? _GEN_31090 : _GEN_28848; // @[rob.scala 166:39]
  wire [6:0] _GEN_33267 = io_i_ex_res_packs_0_valid ? _GEN_31091 : _GEN_28849; // @[rob.scala 166:39]
  wire [6:0] _GEN_33268 = io_i_ex_res_packs_0_valid ? _GEN_31092 : _GEN_28850; // @[rob.scala 166:39]
  wire [6:0] _GEN_33269 = io_i_ex_res_packs_0_valid ? _GEN_31093 : _GEN_28851; // @[rob.scala 166:39]
  wire [6:0] _GEN_33270 = io_i_ex_res_packs_0_valid ? _GEN_31094 : _GEN_28852; // @[rob.scala 166:39]
  wire [6:0] _GEN_33271 = io_i_ex_res_packs_0_valid ? _GEN_31095 : _GEN_28853; // @[rob.scala 166:39]
  wire [6:0] _GEN_33272 = io_i_ex_res_packs_0_valid ? _GEN_31096 : _GEN_28854; // @[rob.scala 166:39]
  wire [6:0] _GEN_33273 = io_i_ex_res_packs_0_valid ? _GEN_31097 : _GEN_28855; // @[rob.scala 166:39]
  wire [6:0] _GEN_33274 = io_i_ex_res_packs_0_valid ? _GEN_31098 : _GEN_28856; // @[rob.scala 166:39]
  wire [6:0] _GEN_33275 = io_i_ex_res_packs_0_valid ? _GEN_31099 : _GEN_28857; // @[rob.scala 166:39]
  wire [6:0] _GEN_33276 = io_i_ex_res_packs_0_valid ? _GEN_31100 : _GEN_28858; // @[rob.scala 166:39]
  wire [6:0] _GEN_33277 = io_i_ex_res_packs_0_valid ? _GEN_31101 : _GEN_28859; // @[rob.scala 166:39]
  wire [6:0] _GEN_33278 = io_i_ex_res_packs_0_valid ? _GEN_31102 : _GEN_28860; // @[rob.scala 166:39]
  wire [6:0] _GEN_33279 = io_i_ex_res_packs_0_valid ? _GEN_31103 : _GEN_28861; // @[rob.scala 166:39]
  wire [6:0] _GEN_33280 = io_i_ex_res_packs_0_valid ? _GEN_31104 : _GEN_28862; // @[rob.scala 166:39]
  wire [6:0] _GEN_33281 = io_i_ex_res_packs_0_valid ? _GEN_31105 : _GEN_28863; // @[rob.scala 166:39]
  wire [6:0] _GEN_33282 = io_i_ex_res_packs_0_valid ? _GEN_31106 : _GEN_28864; // @[rob.scala 166:39]
  wire [6:0] _GEN_33283 = io_i_ex_res_packs_0_valid ? _GEN_31107 : _GEN_28865; // @[rob.scala 166:39]
  wire [6:0] _GEN_33284 = io_i_ex_res_packs_0_valid ? _GEN_31108 : _GEN_28866; // @[rob.scala 166:39]
  wire [6:0] _GEN_33285 = io_i_ex_res_packs_0_valid ? _GEN_31109 : _GEN_28867; // @[rob.scala 166:39]
  wire [6:0] _GEN_33286 = io_i_ex_res_packs_0_valid ? _GEN_31110 : _GEN_28868; // @[rob.scala 166:39]
  wire [6:0] _GEN_33287 = io_i_ex_res_packs_0_valid ? _GEN_31111 : _GEN_28869; // @[rob.scala 166:39]
  wire [6:0] _GEN_33288 = io_i_ex_res_packs_0_valid ? _GEN_31112 : _GEN_28870; // @[rob.scala 166:39]
  wire [6:0] _GEN_33289 = io_i_ex_res_packs_0_valid ? _GEN_31113 : _GEN_28871; // @[rob.scala 166:39]
  wire [6:0] _GEN_33290 = io_i_ex_res_packs_0_valid ? _GEN_31114 : _GEN_28872; // @[rob.scala 166:39]
  wire [6:0] _GEN_33291 = io_i_ex_res_packs_0_valid ? _GEN_31115 : _GEN_28873; // @[rob.scala 166:39]
  wire [6:0] _GEN_33292 = io_i_ex_res_packs_0_valid ? _GEN_31116 : _GEN_28874; // @[rob.scala 166:39]
  wire [6:0] _GEN_33293 = io_i_ex_res_packs_0_valid ? _GEN_31117 : _GEN_28875; // @[rob.scala 166:39]
  wire [6:0] _GEN_33294 = io_i_ex_res_packs_0_valid ? _GEN_31118 : _GEN_28876; // @[rob.scala 166:39]
  wire [6:0] _GEN_33295 = io_i_ex_res_packs_0_valid ? _GEN_31119 : _GEN_28877; // @[rob.scala 166:39]
  wire [6:0] _GEN_33296 = io_i_ex_res_packs_0_valid ? _GEN_31120 : _GEN_28878; // @[rob.scala 166:39]
  wire [6:0] _GEN_33297 = io_i_ex_res_packs_0_valid ? _GEN_31121 : _GEN_28879; // @[rob.scala 166:39]
  wire [6:0] _GEN_33298 = io_i_ex_res_packs_0_valid ? _GEN_31122 : _GEN_28880; // @[rob.scala 166:39]
  wire [6:0] _GEN_33299 = io_i_ex_res_packs_0_valid ? _GEN_31123 : _GEN_28881; // @[rob.scala 166:39]
  wire [6:0] _GEN_33300 = io_i_ex_res_packs_0_valid ? _GEN_31124 : _GEN_28882; // @[rob.scala 166:39]
  wire [6:0] _GEN_33301 = io_i_ex_res_packs_0_valid ? _GEN_31125 : _GEN_28883; // @[rob.scala 166:39]
  wire [6:0] _GEN_33302 = io_i_ex_res_packs_0_valid ? _GEN_31126 : _GEN_28884; // @[rob.scala 166:39]
  wire [6:0] _GEN_33303 = io_i_ex_res_packs_0_valid ? _GEN_31127 : _GEN_28885; // @[rob.scala 166:39]
  wire [6:0] _GEN_33304 = io_i_ex_res_packs_0_valid ? _GEN_31128 : _GEN_28886; // @[rob.scala 166:39]
  wire [6:0] _GEN_33305 = io_i_ex_res_packs_0_valid ? _GEN_31129 : _GEN_28887; // @[rob.scala 166:39]
  wire [6:0] _GEN_33306 = io_i_ex_res_packs_0_valid ? _GEN_31130 : _GEN_28888; // @[rob.scala 166:39]
  wire [6:0] _GEN_33307 = io_i_ex_res_packs_0_valid ? _GEN_31131 : _GEN_28889; // @[rob.scala 166:39]
  wire [6:0] _GEN_33308 = io_i_ex_res_packs_0_valid ? _GEN_31132 : _GEN_28890; // @[rob.scala 166:39]
  wire [6:0] _GEN_33309 = io_i_ex_res_packs_0_valid ? _GEN_31133 : _GEN_28891; // @[rob.scala 166:39]
  wire [6:0] _GEN_33310 = io_i_ex_res_packs_0_valid ? _GEN_31134 : _GEN_28892; // @[rob.scala 166:39]
  wire [6:0] _GEN_33311 = io_i_ex_res_packs_0_valid ? _GEN_31135 : _GEN_28893; // @[rob.scala 166:39]
  wire [6:0] _GEN_33312 = io_i_ex_res_packs_0_valid ? _GEN_31136 : _GEN_28894; // @[rob.scala 166:39]
  wire [6:0] _GEN_33313 = io_i_ex_res_packs_0_valid ? _GEN_31137 : _GEN_28895; // @[rob.scala 166:39]
  wire [6:0] _GEN_33314 = io_i_ex_res_packs_0_valid ? _GEN_31138 : _GEN_28896; // @[rob.scala 166:39]
  wire [6:0] _GEN_33315 = io_i_ex_res_packs_0_valid ? _GEN_31139 : _GEN_28897; // @[rob.scala 166:39]
  wire [6:0] _GEN_33316 = io_i_ex_res_packs_0_valid ? _GEN_31140 : _GEN_28898; // @[rob.scala 166:39]
  wire [6:0] _GEN_33317 = io_i_ex_res_packs_0_valid ? _GEN_31141 : _GEN_28899; // @[rob.scala 166:39]
  wire [6:0] _GEN_33318 = io_i_ex_res_packs_0_valid ? _GEN_31142 : _GEN_28900; // @[rob.scala 166:39]
  wire [6:0] _GEN_33319 = io_i_ex_res_packs_0_valid ? _GEN_31143 : _GEN_28901; // @[rob.scala 166:39]
  wire [6:0] _GEN_33320 = io_i_ex_res_packs_0_valid ? _GEN_31144 : _GEN_28902; // @[rob.scala 166:39]
  wire [6:0] _GEN_33321 = io_i_ex_res_packs_0_valid ? _GEN_31145 : _GEN_28903; // @[rob.scala 166:39]
  wire [6:0] _GEN_33322 = io_i_ex_res_packs_0_valid ? _GEN_31146 : _GEN_28904; // @[rob.scala 166:39]
  wire [6:0] _GEN_33323 = io_i_ex_res_packs_0_valid ? _GEN_31147 : _GEN_28905; // @[rob.scala 166:39]
  wire [6:0] _GEN_33324 = io_i_ex_res_packs_0_valid ? _GEN_31148 : _GEN_28906; // @[rob.scala 166:39]
  wire [6:0] _GEN_33325 = io_i_ex_res_packs_0_valid ? _GEN_31149 : _GEN_28907; // @[rob.scala 166:39]
  wire [6:0] _GEN_33326 = io_i_ex_res_packs_0_valid ? _GEN_31150 : _GEN_28908; // @[rob.scala 166:39]
  wire [6:0] _GEN_33327 = io_i_ex_res_packs_0_valid ? _GEN_31151 : _GEN_28909; // @[rob.scala 166:39]
  wire [6:0] _GEN_33328 = io_i_ex_res_packs_0_valid ? _GEN_31152 : _GEN_28910; // @[rob.scala 166:39]
  wire [6:0] _GEN_33329 = io_i_ex_res_packs_0_valid ? _GEN_31153 : _GEN_28911; // @[rob.scala 166:39]
  wire [6:0] _GEN_33330 = io_i_ex_res_packs_0_valid ? _GEN_31154 : _GEN_28912; // @[rob.scala 166:39]
  wire [6:0] _GEN_33331 = io_i_ex_res_packs_0_valid ? _GEN_31155 : _GEN_28913; // @[rob.scala 166:39]
  wire [6:0] _GEN_33332 = io_i_ex_res_packs_0_valid ? _GEN_31156 : _GEN_28914; // @[rob.scala 166:39]
  wire [6:0] _GEN_33333 = io_i_ex_res_packs_0_valid ? _GEN_31157 : _GEN_28915; // @[rob.scala 166:39]
  wire [6:0] _GEN_33334 = io_i_ex_res_packs_0_valid ? _GEN_31158 : _GEN_28916; // @[rob.scala 166:39]
  wire [6:0] _GEN_33335 = io_i_ex_res_packs_0_valid ? _GEN_31159 : _GEN_28917; // @[rob.scala 166:39]
  wire [6:0] _GEN_33336 = io_i_ex_res_packs_0_valid ? _GEN_31160 : _GEN_28918; // @[rob.scala 166:39]
  wire [6:0] _GEN_33337 = io_i_ex_res_packs_0_valid ? _GEN_31161 : _GEN_28919; // @[rob.scala 166:39]
  wire [6:0] _GEN_33338 = io_i_ex_res_packs_0_valid ? _GEN_31162 : _GEN_28920; // @[rob.scala 166:39]
  wire [6:0] _GEN_33339 = io_i_ex_res_packs_0_valid ? _GEN_31163 : _GEN_28921; // @[rob.scala 166:39]
  wire [6:0] _GEN_33340 = io_i_ex_res_packs_0_valid ? _GEN_31164 : _GEN_28922; // @[rob.scala 166:39]
  wire [6:0] _GEN_33341 = io_i_ex_res_packs_0_valid ? _GEN_31165 : _GEN_28923; // @[rob.scala 166:39]
  wire [6:0] _GEN_33342 = io_i_ex_res_packs_0_valid ? _GEN_31166 : _GEN_28924; // @[rob.scala 166:39]
  wire [6:0] _GEN_33343 = io_i_ex_res_packs_0_valid ? _GEN_31167 : _GEN_28925; // @[rob.scala 166:39]
  wire [6:0] _GEN_33344 = io_i_ex_res_packs_0_valid ? _GEN_31168 : _GEN_28926; // @[rob.scala 166:39]
  wire [6:0] _GEN_33345 = io_i_ex_res_packs_0_valid ? _GEN_31169 : _GEN_28927; // @[rob.scala 166:39]
  wire [6:0] _GEN_33346 = io_i_ex_res_packs_0_valid ? _GEN_31170 : _GEN_28928; // @[rob.scala 166:39]
  wire [6:0] _GEN_33347 = io_i_ex_res_packs_0_valid ? _GEN_31171 : _GEN_28929; // @[rob.scala 166:39]
  wire [6:0] _GEN_33348 = io_i_ex_res_packs_0_valid ? _GEN_31172 : _GEN_28930; // @[rob.scala 166:39]
  wire [6:0] _GEN_33349 = io_i_ex_res_packs_0_valid ? _GEN_31173 : _GEN_28931; // @[rob.scala 166:39]
  wire [4:0] _GEN_33350 = io_i_ex_res_packs_0_valid ? _GEN_31174 : _GEN_28932; // @[rob.scala 166:39]
  wire [4:0] _GEN_33351 = io_i_ex_res_packs_0_valid ? _GEN_31175 : _GEN_28933; // @[rob.scala 166:39]
  wire [4:0] _GEN_33352 = io_i_ex_res_packs_0_valid ? _GEN_31176 : _GEN_28934; // @[rob.scala 166:39]
  wire [4:0] _GEN_33353 = io_i_ex_res_packs_0_valid ? _GEN_31177 : _GEN_28935; // @[rob.scala 166:39]
  wire [4:0] _GEN_33354 = io_i_ex_res_packs_0_valid ? _GEN_31178 : _GEN_28936; // @[rob.scala 166:39]
  wire [4:0] _GEN_33355 = io_i_ex_res_packs_0_valid ? _GEN_31179 : _GEN_28937; // @[rob.scala 166:39]
  wire [4:0] _GEN_33356 = io_i_ex_res_packs_0_valid ? _GEN_31180 : _GEN_28938; // @[rob.scala 166:39]
  wire [4:0] _GEN_33357 = io_i_ex_res_packs_0_valid ? _GEN_31181 : _GEN_28939; // @[rob.scala 166:39]
  wire [4:0] _GEN_33358 = io_i_ex_res_packs_0_valid ? _GEN_31182 : _GEN_28940; // @[rob.scala 166:39]
  wire [4:0] _GEN_33359 = io_i_ex_res_packs_0_valid ? _GEN_31183 : _GEN_28941; // @[rob.scala 166:39]
  wire [4:0] _GEN_33360 = io_i_ex_res_packs_0_valid ? _GEN_31184 : _GEN_28942; // @[rob.scala 166:39]
  wire [4:0] _GEN_33361 = io_i_ex_res_packs_0_valid ? _GEN_31185 : _GEN_28943; // @[rob.scala 166:39]
  wire [4:0] _GEN_33362 = io_i_ex_res_packs_0_valid ? _GEN_31186 : _GEN_28944; // @[rob.scala 166:39]
  wire [4:0] _GEN_33363 = io_i_ex_res_packs_0_valid ? _GEN_31187 : _GEN_28945; // @[rob.scala 166:39]
  wire [4:0] _GEN_33364 = io_i_ex_res_packs_0_valid ? _GEN_31188 : _GEN_28946; // @[rob.scala 166:39]
  wire [4:0] _GEN_33365 = io_i_ex_res_packs_0_valid ? _GEN_31189 : _GEN_28947; // @[rob.scala 166:39]
  wire [4:0] _GEN_33366 = io_i_ex_res_packs_0_valid ? _GEN_31190 : _GEN_28948; // @[rob.scala 166:39]
  wire [4:0] _GEN_33367 = io_i_ex_res_packs_0_valid ? _GEN_31191 : _GEN_28949; // @[rob.scala 166:39]
  wire [4:0] _GEN_33368 = io_i_ex_res_packs_0_valid ? _GEN_31192 : _GEN_28950; // @[rob.scala 166:39]
  wire [4:0] _GEN_33369 = io_i_ex_res_packs_0_valid ? _GEN_31193 : _GEN_28951; // @[rob.scala 166:39]
  wire [4:0] _GEN_33370 = io_i_ex_res_packs_0_valid ? _GEN_31194 : _GEN_28952; // @[rob.scala 166:39]
  wire [4:0] _GEN_33371 = io_i_ex_res_packs_0_valid ? _GEN_31195 : _GEN_28953; // @[rob.scala 166:39]
  wire [4:0] _GEN_33372 = io_i_ex_res_packs_0_valid ? _GEN_31196 : _GEN_28954; // @[rob.scala 166:39]
  wire [4:0] _GEN_33373 = io_i_ex_res_packs_0_valid ? _GEN_31197 : _GEN_28955; // @[rob.scala 166:39]
  wire [4:0] _GEN_33374 = io_i_ex_res_packs_0_valid ? _GEN_31198 : _GEN_28956; // @[rob.scala 166:39]
  wire [4:0] _GEN_33375 = io_i_ex_res_packs_0_valid ? _GEN_31199 : _GEN_28957; // @[rob.scala 166:39]
  wire [4:0] _GEN_33376 = io_i_ex_res_packs_0_valid ? _GEN_31200 : _GEN_28958; // @[rob.scala 166:39]
  wire [4:0] _GEN_33377 = io_i_ex_res_packs_0_valid ? _GEN_31201 : _GEN_28959; // @[rob.scala 166:39]
  wire [4:0] _GEN_33378 = io_i_ex_res_packs_0_valid ? _GEN_31202 : _GEN_28960; // @[rob.scala 166:39]
  wire [4:0] _GEN_33379 = io_i_ex_res_packs_0_valid ? _GEN_31203 : _GEN_28961; // @[rob.scala 166:39]
  wire [4:0] _GEN_33380 = io_i_ex_res_packs_0_valid ? _GEN_31204 : _GEN_28962; // @[rob.scala 166:39]
  wire [4:0] _GEN_33381 = io_i_ex_res_packs_0_valid ? _GEN_31205 : _GEN_28963; // @[rob.scala 166:39]
  wire [4:0] _GEN_33382 = io_i_ex_res_packs_0_valid ? _GEN_31206 : _GEN_28964; // @[rob.scala 166:39]
  wire [4:0] _GEN_33383 = io_i_ex_res_packs_0_valid ? _GEN_31207 : _GEN_28965; // @[rob.scala 166:39]
  wire [4:0] _GEN_33384 = io_i_ex_res_packs_0_valid ? _GEN_31208 : _GEN_28966; // @[rob.scala 166:39]
  wire [4:0] _GEN_33385 = io_i_ex_res_packs_0_valid ? _GEN_31209 : _GEN_28967; // @[rob.scala 166:39]
  wire [4:0] _GEN_33386 = io_i_ex_res_packs_0_valid ? _GEN_31210 : _GEN_28968; // @[rob.scala 166:39]
  wire [4:0] _GEN_33387 = io_i_ex_res_packs_0_valid ? _GEN_31211 : _GEN_28969; // @[rob.scala 166:39]
  wire [4:0] _GEN_33388 = io_i_ex_res_packs_0_valid ? _GEN_31212 : _GEN_28970; // @[rob.scala 166:39]
  wire [4:0] _GEN_33389 = io_i_ex_res_packs_0_valid ? _GEN_31213 : _GEN_28971; // @[rob.scala 166:39]
  wire [4:0] _GEN_33390 = io_i_ex_res_packs_0_valid ? _GEN_31214 : _GEN_28972; // @[rob.scala 166:39]
  wire [4:0] _GEN_33391 = io_i_ex_res_packs_0_valid ? _GEN_31215 : _GEN_28973; // @[rob.scala 166:39]
  wire [4:0] _GEN_33392 = io_i_ex_res_packs_0_valid ? _GEN_31216 : _GEN_28974; // @[rob.scala 166:39]
  wire [4:0] _GEN_33393 = io_i_ex_res_packs_0_valid ? _GEN_31217 : _GEN_28975; // @[rob.scala 166:39]
  wire [4:0] _GEN_33394 = io_i_ex_res_packs_0_valid ? _GEN_31218 : _GEN_28976; // @[rob.scala 166:39]
  wire [4:0] _GEN_33395 = io_i_ex_res_packs_0_valid ? _GEN_31219 : _GEN_28977; // @[rob.scala 166:39]
  wire [4:0] _GEN_33396 = io_i_ex_res_packs_0_valid ? _GEN_31220 : _GEN_28978; // @[rob.scala 166:39]
  wire [4:0] _GEN_33397 = io_i_ex_res_packs_0_valid ? _GEN_31221 : _GEN_28979; // @[rob.scala 166:39]
  wire [4:0] _GEN_33398 = io_i_ex_res_packs_0_valid ? _GEN_31222 : _GEN_28980; // @[rob.scala 166:39]
  wire [4:0] _GEN_33399 = io_i_ex_res_packs_0_valid ? _GEN_31223 : _GEN_28981; // @[rob.scala 166:39]
  wire [4:0] _GEN_33400 = io_i_ex_res_packs_0_valid ? _GEN_31224 : _GEN_28982; // @[rob.scala 166:39]
  wire [4:0] _GEN_33401 = io_i_ex_res_packs_0_valid ? _GEN_31225 : _GEN_28983; // @[rob.scala 166:39]
  wire [4:0] _GEN_33402 = io_i_ex_res_packs_0_valid ? _GEN_31226 : _GEN_28984; // @[rob.scala 166:39]
  wire [4:0] _GEN_33403 = io_i_ex_res_packs_0_valid ? _GEN_31227 : _GEN_28985; // @[rob.scala 166:39]
  wire [4:0] _GEN_33404 = io_i_ex_res_packs_0_valid ? _GEN_31228 : _GEN_28986; // @[rob.scala 166:39]
  wire [4:0] _GEN_33405 = io_i_ex_res_packs_0_valid ? _GEN_31229 : _GEN_28987; // @[rob.scala 166:39]
  wire [4:0] _GEN_33406 = io_i_ex_res_packs_0_valid ? _GEN_31230 : _GEN_28988; // @[rob.scala 166:39]
  wire [4:0] _GEN_33407 = io_i_ex_res_packs_0_valid ? _GEN_31231 : _GEN_28989; // @[rob.scala 166:39]
  wire [4:0] _GEN_33408 = io_i_ex_res_packs_0_valid ? _GEN_31232 : _GEN_28990; // @[rob.scala 166:39]
  wire [4:0] _GEN_33409 = io_i_ex_res_packs_0_valid ? _GEN_31233 : _GEN_28991; // @[rob.scala 166:39]
  wire [4:0] _GEN_33410 = io_i_ex_res_packs_0_valid ? _GEN_31234 : _GEN_28992; // @[rob.scala 166:39]
  wire [4:0] _GEN_33411 = io_i_ex_res_packs_0_valid ? _GEN_31235 : _GEN_28993; // @[rob.scala 166:39]
  wire [4:0] _GEN_33412 = io_i_ex_res_packs_0_valid ? _GEN_31236 : _GEN_28994; // @[rob.scala 166:39]
  wire [4:0] _GEN_33413 = io_i_ex_res_packs_0_valid ? _GEN_31237 : _GEN_28995; // @[rob.scala 166:39]
  wire [63:0] _GEN_34054 = io_i_ex_res_packs_0_valid ? _GEN_31878 : _GEN_29636; // @[rob.scala 166:39]
  wire [63:0] _GEN_34055 = io_i_ex_res_packs_0_valid ? _GEN_31879 : _GEN_29637; // @[rob.scala 166:39]
  wire [63:0] _GEN_34056 = io_i_ex_res_packs_0_valid ? _GEN_31880 : _GEN_29638; // @[rob.scala 166:39]
  wire [63:0] _GEN_34057 = io_i_ex_res_packs_0_valid ? _GEN_31881 : _GEN_29639; // @[rob.scala 166:39]
  wire [63:0] _GEN_34058 = io_i_ex_res_packs_0_valid ? _GEN_31882 : _GEN_29640; // @[rob.scala 166:39]
  wire [63:0] _GEN_34059 = io_i_ex_res_packs_0_valid ? _GEN_31883 : _GEN_29641; // @[rob.scala 166:39]
  wire [63:0] _GEN_34060 = io_i_ex_res_packs_0_valid ? _GEN_31884 : _GEN_29642; // @[rob.scala 166:39]
  wire [63:0] _GEN_34061 = io_i_ex_res_packs_0_valid ? _GEN_31885 : _GEN_29643; // @[rob.scala 166:39]
  wire [63:0] _GEN_34062 = io_i_ex_res_packs_0_valid ? _GEN_31886 : _GEN_29644; // @[rob.scala 166:39]
  wire [63:0] _GEN_34063 = io_i_ex_res_packs_0_valid ? _GEN_31887 : _GEN_29645; // @[rob.scala 166:39]
  wire [63:0] _GEN_34064 = io_i_ex_res_packs_0_valid ? _GEN_31888 : _GEN_29646; // @[rob.scala 166:39]
  wire [63:0] _GEN_34065 = io_i_ex_res_packs_0_valid ? _GEN_31889 : _GEN_29647; // @[rob.scala 166:39]
  wire [63:0] _GEN_34066 = io_i_ex_res_packs_0_valid ? _GEN_31890 : _GEN_29648; // @[rob.scala 166:39]
  wire [63:0] _GEN_34067 = io_i_ex_res_packs_0_valid ? _GEN_31891 : _GEN_29649; // @[rob.scala 166:39]
  wire [63:0] _GEN_34068 = io_i_ex_res_packs_0_valid ? _GEN_31892 : _GEN_29650; // @[rob.scala 166:39]
  wire [63:0] _GEN_34069 = io_i_ex_res_packs_0_valid ? _GEN_31893 : _GEN_29651; // @[rob.scala 166:39]
  wire [63:0] _GEN_34070 = io_i_ex_res_packs_0_valid ? _GEN_31894 : _GEN_29652; // @[rob.scala 166:39]
  wire [63:0] _GEN_34071 = io_i_ex_res_packs_0_valid ? _GEN_31895 : _GEN_29653; // @[rob.scala 166:39]
  wire [63:0] _GEN_34072 = io_i_ex_res_packs_0_valid ? _GEN_31896 : _GEN_29654; // @[rob.scala 166:39]
  wire [63:0] _GEN_34073 = io_i_ex_res_packs_0_valid ? _GEN_31897 : _GEN_29655; // @[rob.scala 166:39]
  wire [63:0] _GEN_34074 = io_i_ex_res_packs_0_valid ? _GEN_31898 : _GEN_29656; // @[rob.scala 166:39]
  wire [63:0] _GEN_34075 = io_i_ex_res_packs_0_valid ? _GEN_31899 : _GEN_29657; // @[rob.scala 166:39]
  wire [63:0] _GEN_34076 = io_i_ex_res_packs_0_valid ? _GEN_31900 : _GEN_29658; // @[rob.scala 166:39]
  wire [63:0] _GEN_34077 = io_i_ex_res_packs_0_valid ? _GEN_31901 : _GEN_29659; // @[rob.scala 166:39]
  wire [63:0] _GEN_34078 = io_i_ex_res_packs_0_valid ? _GEN_31902 : _GEN_29660; // @[rob.scala 166:39]
  wire [63:0] _GEN_34079 = io_i_ex_res_packs_0_valid ? _GEN_31903 : _GEN_29661; // @[rob.scala 166:39]
  wire [63:0] _GEN_34080 = io_i_ex_res_packs_0_valid ? _GEN_31904 : _GEN_29662; // @[rob.scala 166:39]
  wire [63:0] _GEN_34081 = io_i_ex_res_packs_0_valid ? _GEN_31905 : _GEN_29663; // @[rob.scala 166:39]
  wire [63:0] _GEN_34082 = io_i_ex_res_packs_0_valid ? _GEN_31906 : _GEN_29664; // @[rob.scala 166:39]
  wire [63:0] _GEN_34083 = io_i_ex_res_packs_0_valid ? _GEN_31907 : _GEN_29665; // @[rob.scala 166:39]
  wire [63:0] _GEN_34084 = io_i_ex_res_packs_0_valid ? _GEN_31908 : _GEN_29666; // @[rob.scala 166:39]
  wire [63:0] _GEN_34085 = io_i_ex_res_packs_0_valid ? _GEN_31909 : _GEN_29667; // @[rob.scala 166:39]
  wire [63:0] _GEN_34086 = io_i_ex_res_packs_0_valid ? _GEN_31910 : _GEN_29668; // @[rob.scala 166:39]
  wire [63:0] _GEN_34087 = io_i_ex_res_packs_0_valid ? _GEN_31911 : _GEN_29669; // @[rob.scala 166:39]
  wire [63:0] _GEN_34088 = io_i_ex_res_packs_0_valid ? _GEN_31912 : _GEN_29670; // @[rob.scala 166:39]
  wire [63:0] _GEN_34089 = io_i_ex_res_packs_0_valid ? _GEN_31913 : _GEN_29671; // @[rob.scala 166:39]
  wire [63:0] _GEN_34090 = io_i_ex_res_packs_0_valid ? _GEN_31914 : _GEN_29672; // @[rob.scala 166:39]
  wire [63:0] _GEN_34091 = io_i_ex_res_packs_0_valid ? _GEN_31915 : _GEN_29673; // @[rob.scala 166:39]
  wire [63:0] _GEN_34092 = io_i_ex_res_packs_0_valid ? _GEN_31916 : _GEN_29674; // @[rob.scala 166:39]
  wire [63:0] _GEN_34093 = io_i_ex_res_packs_0_valid ? _GEN_31917 : _GEN_29675; // @[rob.scala 166:39]
  wire [63:0] _GEN_34094 = io_i_ex_res_packs_0_valid ? _GEN_31918 : _GEN_29676; // @[rob.scala 166:39]
  wire [63:0] _GEN_34095 = io_i_ex_res_packs_0_valid ? _GEN_31919 : _GEN_29677; // @[rob.scala 166:39]
  wire [63:0] _GEN_34096 = io_i_ex_res_packs_0_valid ? _GEN_31920 : _GEN_29678; // @[rob.scala 166:39]
  wire [63:0] _GEN_34097 = io_i_ex_res_packs_0_valid ? _GEN_31921 : _GEN_29679; // @[rob.scala 166:39]
  wire [63:0] _GEN_34098 = io_i_ex_res_packs_0_valid ? _GEN_31922 : _GEN_29680; // @[rob.scala 166:39]
  wire [63:0] _GEN_34099 = io_i_ex_res_packs_0_valid ? _GEN_31923 : _GEN_29681; // @[rob.scala 166:39]
  wire [63:0] _GEN_34100 = io_i_ex_res_packs_0_valid ? _GEN_31924 : _GEN_29682; // @[rob.scala 166:39]
  wire [63:0] _GEN_34101 = io_i_ex_res_packs_0_valid ? _GEN_31925 : _GEN_29683; // @[rob.scala 166:39]
  wire [63:0] _GEN_34102 = io_i_ex_res_packs_0_valid ? _GEN_31926 : _GEN_29684; // @[rob.scala 166:39]
  wire [63:0] _GEN_34103 = io_i_ex_res_packs_0_valid ? _GEN_31927 : _GEN_29685; // @[rob.scala 166:39]
  wire [63:0] _GEN_34104 = io_i_ex_res_packs_0_valid ? _GEN_31928 : _GEN_29686; // @[rob.scala 166:39]
  wire [63:0] _GEN_34105 = io_i_ex_res_packs_0_valid ? _GEN_31929 : _GEN_29687; // @[rob.scala 166:39]
  wire [63:0] _GEN_34106 = io_i_ex_res_packs_0_valid ? _GEN_31930 : _GEN_29688; // @[rob.scala 166:39]
  wire [63:0] _GEN_34107 = io_i_ex_res_packs_0_valid ? _GEN_31931 : _GEN_29689; // @[rob.scala 166:39]
  wire [63:0] _GEN_34108 = io_i_ex_res_packs_0_valid ? _GEN_31932 : _GEN_29690; // @[rob.scala 166:39]
  wire [63:0] _GEN_34109 = io_i_ex_res_packs_0_valid ? _GEN_31933 : _GEN_29691; // @[rob.scala 166:39]
  wire [63:0] _GEN_34110 = io_i_ex_res_packs_0_valid ? _GEN_31934 : _GEN_29692; // @[rob.scala 166:39]
  wire [63:0] _GEN_34111 = io_i_ex_res_packs_0_valid ? _GEN_31935 : _GEN_29693; // @[rob.scala 166:39]
  wire [63:0] _GEN_34112 = io_i_ex_res_packs_0_valid ? _GEN_31936 : _GEN_29694; // @[rob.scala 166:39]
  wire [63:0] _GEN_34113 = io_i_ex_res_packs_0_valid ? _GEN_31937 : _GEN_29695; // @[rob.scala 166:39]
  wire [63:0] _GEN_34114 = io_i_ex_res_packs_0_valid ? _GEN_31938 : _GEN_29696; // @[rob.scala 166:39]
  wire [63:0] _GEN_34115 = io_i_ex_res_packs_0_valid ? _GEN_31939 : _GEN_29697; // @[rob.scala 166:39]
  wire [63:0] _GEN_34116 = io_i_ex_res_packs_0_valid ? _GEN_31940 : _GEN_29698; // @[rob.scala 166:39]
  wire [63:0] _GEN_34117 = io_i_ex_res_packs_0_valid ? _GEN_31941 : _GEN_29699; // @[rob.scala 166:39]
  wire [63:0] _GEN_34118 = io_i_ex_res_packs_0_valid ? _GEN_31942 : _GEN_29700; // @[rob.scala 166:39]
  wire [63:0] _GEN_34119 = io_i_ex_res_packs_0_valid ? _GEN_31943 : _GEN_29701; // @[rob.scala 166:39]
  wire [63:0] _GEN_34120 = io_i_ex_res_packs_0_valid ? _GEN_31944 : _GEN_29702; // @[rob.scala 166:39]
  wire [63:0] _GEN_34121 = io_i_ex_res_packs_0_valid ? _GEN_31945 : _GEN_29703; // @[rob.scala 166:39]
  wire [63:0] _GEN_34122 = io_i_ex_res_packs_0_valid ? _GEN_31946 : _GEN_29704; // @[rob.scala 166:39]
  wire [63:0] _GEN_34123 = io_i_ex_res_packs_0_valid ? _GEN_31947 : _GEN_29705; // @[rob.scala 166:39]
  wire [63:0] _GEN_34124 = io_i_ex_res_packs_0_valid ? _GEN_31948 : _GEN_29706; // @[rob.scala 166:39]
  wire [63:0] _GEN_34125 = io_i_ex_res_packs_0_valid ? _GEN_31949 : _GEN_29707; // @[rob.scala 166:39]
  wire [63:0] _GEN_34126 = io_i_ex_res_packs_0_valid ? _GEN_31950 : _GEN_29708; // @[rob.scala 166:39]
  wire [63:0] _GEN_34127 = io_i_ex_res_packs_0_valid ? _GEN_31951 : _GEN_29709; // @[rob.scala 166:39]
  wire [63:0] _GEN_34128 = io_i_ex_res_packs_0_valid ? _GEN_31952 : _GEN_29710; // @[rob.scala 166:39]
  wire [63:0] _GEN_34129 = io_i_ex_res_packs_0_valid ? _GEN_31953 : _GEN_29711; // @[rob.scala 166:39]
  wire [63:0] _GEN_34130 = io_i_ex_res_packs_0_valid ? _GEN_31954 : _GEN_29712; // @[rob.scala 166:39]
  wire [63:0] _GEN_34131 = io_i_ex_res_packs_0_valid ? _GEN_31955 : _GEN_29713; // @[rob.scala 166:39]
  wire [63:0] _GEN_34132 = io_i_ex_res_packs_0_valid ? _GEN_31956 : _GEN_29714; // @[rob.scala 166:39]
  wire [63:0] _GEN_34133 = io_i_ex_res_packs_0_valid ? _GEN_31957 : _GEN_29715; // @[rob.scala 166:39]
  wire [63:0] _GEN_34134 = io_i_ex_res_packs_0_valid ? _GEN_31958 : _GEN_29716; // @[rob.scala 166:39]
  wire [63:0] _GEN_34135 = io_i_ex_res_packs_0_valid ? _GEN_31959 : _GEN_29717; // @[rob.scala 166:39]
  wire [63:0] _GEN_34136 = io_i_ex_res_packs_0_valid ? _GEN_31960 : _GEN_29718; // @[rob.scala 166:39]
  wire [63:0] _GEN_34137 = io_i_ex_res_packs_0_valid ? _GEN_31961 : _GEN_29719; // @[rob.scala 166:39]
  wire [63:0] _GEN_34138 = io_i_ex_res_packs_0_valid ? _GEN_31962 : _GEN_29720; // @[rob.scala 166:39]
  wire [63:0] _GEN_34139 = io_i_ex_res_packs_0_valid ? _GEN_31963 : _GEN_29721; // @[rob.scala 166:39]
  wire [63:0] _GEN_34140 = io_i_ex_res_packs_0_valid ? _GEN_31964 : _GEN_29722; // @[rob.scala 166:39]
  wire [63:0] _GEN_34141 = io_i_ex_res_packs_0_valid ? _GEN_31965 : _GEN_29723; // @[rob.scala 166:39]
  wire [63:0] _GEN_34142 = io_i_ex_res_packs_0_valid ? _GEN_31966 : _GEN_29724; // @[rob.scala 166:39]
  wire [63:0] _GEN_34143 = io_i_ex_res_packs_0_valid ? _GEN_31967 : _GEN_29725; // @[rob.scala 166:39]
  wire [63:0] _GEN_34144 = io_i_ex_res_packs_0_valid ? _GEN_31968 : _GEN_29726; // @[rob.scala 166:39]
  wire [63:0] _GEN_34145 = io_i_ex_res_packs_0_valid ? _GEN_31969 : _GEN_29727; // @[rob.scala 166:39]
  wire [63:0] _GEN_34146 = io_i_ex_res_packs_0_valid ? _GEN_31970 : _GEN_29728; // @[rob.scala 166:39]
  wire [63:0] _GEN_34147 = io_i_ex_res_packs_0_valid ? _GEN_31971 : _GEN_29729; // @[rob.scala 166:39]
  wire [63:0] _GEN_34148 = io_i_ex_res_packs_0_valid ? _GEN_31972 : _GEN_29730; // @[rob.scala 166:39]
  wire [63:0] _GEN_34149 = io_i_ex_res_packs_0_valid ? _GEN_31973 : _GEN_29731; // @[rob.scala 166:39]
  wire [63:0] _GEN_34150 = io_i_ex_res_packs_0_valid ? _GEN_31974 : _GEN_29732; // @[rob.scala 166:39]
  wire [63:0] _GEN_34151 = io_i_ex_res_packs_0_valid ? _GEN_31975 : _GEN_29733; // @[rob.scala 166:39]
  wire [63:0] _GEN_34152 = io_i_ex_res_packs_0_valid ? _GEN_31976 : _GEN_29734; // @[rob.scala 166:39]
  wire [63:0] _GEN_34153 = io_i_ex_res_packs_0_valid ? _GEN_31977 : _GEN_29735; // @[rob.scala 166:39]
  wire [63:0] _GEN_34154 = io_i_ex_res_packs_0_valid ? _GEN_31978 : _GEN_29736; // @[rob.scala 166:39]
  wire [63:0] _GEN_34155 = io_i_ex_res_packs_0_valid ? _GEN_31979 : _GEN_29737; // @[rob.scala 166:39]
  wire [63:0] _GEN_34156 = io_i_ex_res_packs_0_valid ? _GEN_31980 : _GEN_29738; // @[rob.scala 166:39]
  wire [63:0] _GEN_34157 = io_i_ex_res_packs_0_valid ? _GEN_31981 : _GEN_29739; // @[rob.scala 166:39]
  wire [63:0] _GEN_34158 = io_i_ex_res_packs_0_valid ? _GEN_31982 : _GEN_29740; // @[rob.scala 166:39]
  wire [63:0] _GEN_34159 = io_i_ex_res_packs_0_valid ? _GEN_31983 : _GEN_29741; // @[rob.scala 166:39]
  wire [63:0] _GEN_34160 = io_i_ex_res_packs_0_valid ? _GEN_31984 : _GEN_29742; // @[rob.scala 166:39]
  wire [63:0] _GEN_34161 = io_i_ex_res_packs_0_valid ? _GEN_31985 : _GEN_29743; // @[rob.scala 166:39]
  wire [63:0] _GEN_34162 = io_i_ex_res_packs_0_valid ? _GEN_31986 : _GEN_29744; // @[rob.scala 166:39]
  wire [63:0] _GEN_34163 = io_i_ex_res_packs_0_valid ? _GEN_31987 : _GEN_29745; // @[rob.scala 166:39]
  wire [63:0] _GEN_34164 = io_i_ex_res_packs_0_valid ? _GEN_31988 : _GEN_29746; // @[rob.scala 166:39]
  wire [63:0] _GEN_34165 = io_i_ex_res_packs_0_valid ? _GEN_31989 : _GEN_29747; // @[rob.scala 166:39]
  wire [63:0] _GEN_34166 = io_i_ex_res_packs_0_valid ? _GEN_31990 : _GEN_29748; // @[rob.scala 166:39]
  wire [63:0] _GEN_34167 = io_i_ex_res_packs_0_valid ? _GEN_31991 : _GEN_29749; // @[rob.scala 166:39]
  wire [63:0] _GEN_34168 = io_i_ex_res_packs_0_valid ? _GEN_31992 : _GEN_29750; // @[rob.scala 166:39]
  wire [63:0] _GEN_34169 = io_i_ex_res_packs_0_valid ? _GEN_31993 : _GEN_29751; // @[rob.scala 166:39]
  wire [63:0] _GEN_34170 = io_i_ex_res_packs_0_valid ? _GEN_31994 : _GEN_29752; // @[rob.scala 166:39]
  wire [63:0] _GEN_34171 = io_i_ex_res_packs_0_valid ? _GEN_31995 : _GEN_29753; // @[rob.scala 166:39]
  wire [63:0] _GEN_34172 = io_i_ex_res_packs_0_valid ? _GEN_31996 : _GEN_29754; // @[rob.scala 166:39]
  wire [63:0] _GEN_34173 = io_i_ex_res_packs_0_valid ? _GEN_31997 : _GEN_29755; // @[rob.scala 166:39]
  wire [63:0] _GEN_34174 = io_i_ex_res_packs_0_valid ? _GEN_31998 : _GEN_29756; // @[rob.scala 166:39]
  wire [63:0] _GEN_34175 = io_i_ex_res_packs_0_valid ? _GEN_31999 : _GEN_29757; // @[rob.scala 166:39]
  wire [63:0] _GEN_34176 = io_i_ex_res_packs_0_valid ? _GEN_32000 : _GEN_29758; // @[rob.scala 166:39]
  wire [63:0] _GEN_34177 = io_i_ex_res_packs_0_valid ? _GEN_32001 : _GEN_29759; // @[rob.scala 166:39]
  wire [63:0] _GEN_34178 = io_i_ex_res_packs_0_valid ? _GEN_32002 : _GEN_29760; // @[rob.scala 166:39]
  wire [63:0] _GEN_34179 = io_i_ex_res_packs_0_valid ? _GEN_32003 : _GEN_29761; // @[rob.scala 166:39]
  wire [63:0] _GEN_34180 = io_i_ex_res_packs_0_valid ? _GEN_32004 : _GEN_29762; // @[rob.scala 166:39]
  wire [63:0] _GEN_34181 = io_i_ex_res_packs_0_valid ? _GEN_32005 : _GEN_29763; // @[rob.scala 166:39]
  wire [4:0] _GEN_34438 = io_i_ex_res_packs_0_valid ? _GEN_32262 : _GEN_30020; // @[rob.scala 166:39]
  wire [4:0] _GEN_34439 = io_i_ex_res_packs_0_valid ? _GEN_32263 : _GEN_30021; // @[rob.scala 166:39]
  wire [4:0] _GEN_34440 = io_i_ex_res_packs_0_valid ? _GEN_32264 : _GEN_30022; // @[rob.scala 166:39]
  wire [4:0] _GEN_34441 = io_i_ex_res_packs_0_valid ? _GEN_32265 : _GEN_30023; // @[rob.scala 166:39]
  wire [4:0] _GEN_34442 = io_i_ex_res_packs_0_valid ? _GEN_32266 : _GEN_30024; // @[rob.scala 166:39]
  wire [4:0] _GEN_34443 = io_i_ex_res_packs_0_valid ? _GEN_32267 : _GEN_30025; // @[rob.scala 166:39]
  wire [4:0] _GEN_34444 = io_i_ex_res_packs_0_valid ? _GEN_32268 : _GEN_30026; // @[rob.scala 166:39]
  wire [4:0] _GEN_34445 = io_i_ex_res_packs_0_valid ? _GEN_32269 : _GEN_30027; // @[rob.scala 166:39]
  wire [4:0] _GEN_34446 = io_i_ex_res_packs_0_valid ? _GEN_32270 : _GEN_30028; // @[rob.scala 166:39]
  wire [4:0] _GEN_34447 = io_i_ex_res_packs_0_valid ? _GEN_32271 : _GEN_30029; // @[rob.scala 166:39]
  wire [4:0] _GEN_34448 = io_i_ex_res_packs_0_valid ? _GEN_32272 : _GEN_30030; // @[rob.scala 166:39]
  wire [4:0] _GEN_34449 = io_i_ex_res_packs_0_valid ? _GEN_32273 : _GEN_30031; // @[rob.scala 166:39]
  wire [4:0] _GEN_34450 = io_i_ex_res_packs_0_valid ? _GEN_32274 : _GEN_30032; // @[rob.scala 166:39]
  wire [4:0] _GEN_34451 = io_i_ex_res_packs_0_valid ? _GEN_32275 : _GEN_30033; // @[rob.scala 166:39]
  wire [4:0] _GEN_34452 = io_i_ex_res_packs_0_valid ? _GEN_32276 : _GEN_30034; // @[rob.scala 166:39]
  wire [4:0] _GEN_34453 = io_i_ex_res_packs_0_valid ? _GEN_32277 : _GEN_30035; // @[rob.scala 166:39]
  wire [4:0] _GEN_34454 = io_i_ex_res_packs_0_valid ? _GEN_32278 : _GEN_30036; // @[rob.scala 166:39]
  wire [4:0] _GEN_34455 = io_i_ex_res_packs_0_valid ? _GEN_32279 : _GEN_30037; // @[rob.scala 166:39]
  wire [4:0] _GEN_34456 = io_i_ex_res_packs_0_valid ? _GEN_32280 : _GEN_30038; // @[rob.scala 166:39]
  wire [4:0] _GEN_34457 = io_i_ex_res_packs_0_valid ? _GEN_32281 : _GEN_30039; // @[rob.scala 166:39]
  wire [4:0] _GEN_34458 = io_i_ex_res_packs_0_valid ? _GEN_32282 : _GEN_30040; // @[rob.scala 166:39]
  wire [4:0] _GEN_34459 = io_i_ex_res_packs_0_valid ? _GEN_32283 : _GEN_30041; // @[rob.scala 166:39]
  wire [4:0] _GEN_34460 = io_i_ex_res_packs_0_valid ? _GEN_32284 : _GEN_30042; // @[rob.scala 166:39]
  wire [4:0] _GEN_34461 = io_i_ex_res_packs_0_valid ? _GEN_32285 : _GEN_30043; // @[rob.scala 166:39]
  wire [4:0] _GEN_34462 = io_i_ex_res_packs_0_valid ? _GEN_32286 : _GEN_30044; // @[rob.scala 166:39]
  wire [4:0] _GEN_34463 = io_i_ex_res_packs_0_valid ? _GEN_32287 : _GEN_30045; // @[rob.scala 166:39]
  wire [4:0] _GEN_34464 = io_i_ex_res_packs_0_valid ? _GEN_32288 : _GEN_30046; // @[rob.scala 166:39]
  wire [4:0] _GEN_34465 = io_i_ex_res_packs_0_valid ? _GEN_32289 : _GEN_30047; // @[rob.scala 166:39]
  wire [4:0] _GEN_34466 = io_i_ex_res_packs_0_valid ? _GEN_32290 : _GEN_30048; // @[rob.scala 166:39]
  wire [4:0] _GEN_34467 = io_i_ex_res_packs_0_valid ? _GEN_32291 : _GEN_30049; // @[rob.scala 166:39]
  wire [4:0] _GEN_34468 = io_i_ex_res_packs_0_valid ? _GEN_32292 : _GEN_30050; // @[rob.scala 166:39]
  wire [4:0] _GEN_34469 = io_i_ex_res_packs_0_valid ? _GEN_32293 : _GEN_30051; // @[rob.scala 166:39]
  wire [4:0] _GEN_34470 = io_i_ex_res_packs_0_valid ? _GEN_32294 : _GEN_30052; // @[rob.scala 166:39]
  wire [4:0] _GEN_34471 = io_i_ex_res_packs_0_valid ? _GEN_32295 : _GEN_30053; // @[rob.scala 166:39]
  wire [4:0] _GEN_34472 = io_i_ex_res_packs_0_valid ? _GEN_32296 : _GEN_30054; // @[rob.scala 166:39]
  wire [4:0] _GEN_34473 = io_i_ex_res_packs_0_valid ? _GEN_32297 : _GEN_30055; // @[rob.scala 166:39]
  wire [4:0] _GEN_34474 = io_i_ex_res_packs_0_valid ? _GEN_32298 : _GEN_30056; // @[rob.scala 166:39]
  wire [4:0] _GEN_34475 = io_i_ex_res_packs_0_valid ? _GEN_32299 : _GEN_30057; // @[rob.scala 166:39]
  wire [4:0] _GEN_34476 = io_i_ex_res_packs_0_valid ? _GEN_32300 : _GEN_30058; // @[rob.scala 166:39]
  wire [4:0] _GEN_34477 = io_i_ex_res_packs_0_valid ? _GEN_32301 : _GEN_30059; // @[rob.scala 166:39]
  wire [4:0] _GEN_34478 = io_i_ex_res_packs_0_valid ? _GEN_32302 : _GEN_30060; // @[rob.scala 166:39]
  wire [4:0] _GEN_34479 = io_i_ex_res_packs_0_valid ? _GEN_32303 : _GEN_30061; // @[rob.scala 166:39]
  wire [4:0] _GEN_34480 = io_i_ex_res_packs_0_valid ? _GEN_32304 : _GEN_30062; // @[rob.scala 166:39]
  wire [4:0] _GEN_34481 = io_i_ex_res_packs_0_valid ? _GEN_32305 : _GEN_30063; // @[rob.scala 166:39]
  wire [4:0] _GEN_34482 = io_i_ex_res_packs_0_valid ? _GEN_32306 : _GEN_30064; // @[rob.scala 166:39]
  wire [4:0] _GEN_34483 = io_i_ex_res_packs_0_valid ? _GEN_32307 : _GEN_30065; // @[rob.scala 166:39]
  wire [4:0] _GEN_34484 = io_i_ex_res_packs_0_valid ? _GEN_32308 : _GEN_30066; // @[rob.scala 166:39]
  wire [4:0] _GEN_34485 = io_i_ex_res_packs_0_valid ? _GEN_32309 : _GEN_30067; // @[rob.scala 166:39]
  wire [4:0] _GEN_34486 = io_i_ex_res_packs_0_valid ? _GEN_32310 : _GEN_30068; // @[rob.scala 166:39]
  wire [4:0] _GEN_34487 = io_i_ex_res_packs_0_valid ? _GEN_32311 : _GEN_30069; // @[rob.scala 166:39]
  wire [4:0] _GEN_34488 = io_i_ex_res_packs_0_valid ? _GEN_32312 : _GEN_30070; // @[rob.scala 166:39]
  wire [4:0] _GEN_34489 = io_i_ex_res_packs_0_valid ? _GEN_32313 : _GEN_30071; // @[rob.scala 166:39]
  wire [4:0] _GEN_34490 = io_i_ex_res_packs_0_valid ? _GEN_32314 : _GEN_30072; // @[rob.scala 166:39]
  wire [4:0] _GEN_34491 = io_i_ex_res_packs_0_valid ? _GEN_32315 : _GEN_30073; // @[rob.scala 166:39]
  wire [4:0] _GEN_34492 = io_i_ex_res_packs_0_valid ? _GEN_32316 : _GEN_30074; // @[rob.scala 166:39]
  wire [4:0] _GEN_34493 = io_i_ex_res_packs_0_valid ? _GEN_32317 : _GEN_30075; // @[rob.scala 166:39]
  wire [4:0] _GEN_34494 = io_i_ex_res_packs_0_valid ? _GEN_32318 : _GEN_30076; // @[rob.scala 166:39]
  wire [4:0] _GEN_34495 = io_i_ex_res_packs_0_valid ? _GEN_32319 : _GEN_30077; // @[rob.scala 166:39]
  wire [4:0] _GEN_34496 = io_i_ex_res_packs_0_valid ? _GEN_32320 : _GEN_30078; // @[rob.scala 166:39]
  wire [4:0] _GEN_34497 = io_i_ex_res_packs_0_valid ? _GEN_32321 : _GEN_30079; // @[rob.scala 166:39]
  wire [4:0] _GEN_34498 = io_i_ex_res_packs_0_valid ? _GEN_32322 : _GEN_30080; // @[rob.scala 166:39]
  wire [4:0] _GEN_34499 = io_i_ex_res_packs_0_valid ? _GEN_32323 : _GEN_30081; // @[rob.scala 166:39]
  wire [4:0] _GEN_34500 = io_i_ex_res_packs_0_valid ? _GEN_32324 : _GEN_30082; // @[rob.scala 166:39]
  wire [4:0] _GEN_34501 = io_i_ex_res_packs_0_valid ? _GEN_32325 : _GEN_30083; // @[rob.scala 166:39]
  wire  _GEN_34694 = io_i_ex_res_packs_0_valid ? _GEN_32518 : _GEN_30276; // @[rob.scala 166:39]
  wire  _GEN_34695 = io_i_ex_res_packs_0_valid ? _GEN_32519 : _GEN_30277; // @[rob.scala 166:39]
  wire  _GEN_34696 = io_i_ex_res_packs_0_valid ? _GEN_32520 : _GEN_30278; // @[rob.scala 166:39]
  wire  _GEN_34697 = io_i_ex_res_packs_0_valid ? _GEN_32521 : _GEN_30279; // @[rob.scala 166:39]
  wire  _GEN_34698 = io_i_ex_res_packs_0_valid ? _GEN_32522 : _GEN_30280; // @[rob.scala 166:39]
  wire  _GEN_34699 = io_i_ex_res_packs_0_valid ? _GEN_32523 : _GEN_30281; // @[rob.scala 166:39]
  wire  _GEN_34700 = io_i_ex_res_packs_0_valid ? _GEN_32524 : _GEN_30282; // @[rob.scala 166:39]
  wire  _GEN_34701 = io_i_ex_res_packs_0_valid ? _GEN_32525 : _GEN_30283; // @[rob.scala 166:39]
  wire  _GEN_34702 = io_i_ex_res_packs_0_valid ? _GEN_32526 : _GEN_30284; // @[rob.scala 166:39]
  wire  _GEN_34703 = io_i_ex_res_packs_0_valid ? _GEN_32527 : _GEN_30285; // @[rob.scala 166:39]
  wire  _GEN_34704 = io_i_ex_res_packs_0_valid ? _GEN_32528 : _GEN_30286; // @[rob.scala 166:39]
  wire  _GEN_34705 = io_i_ex_res_packs_0_valid ? _GEN_32529 : _GEN_30287; // @[rob.scala 166:39]
  wire  _GEN_34706 = io_i_ex_res_packs_0_valid ? _GEN_32530 : _GEN_30288; // @[rob.scala 166:39]
  wire  _GEN_34707 = io_i_ex_res_packs_0_valid ? _GEN_32531 : _GEN_30289; // @[rob.scala 166:39]
  wire  _GEN_34708 = io_i_ex_res_packs_0_valid ? _GEN_32532 : _GEN_30290; // @[rob.scala 166:39]
  wire  _GEN_34709 = io_i_ex_res_packs_0_valid ? _GEN_32533 : _GEN_30291; // @[rob.scala 166:39]
  wire  _GEN_34710 = io_i_ex_res_packs_0_valid ? _GEN_32534 : _GEN_30292; // @[rob.scala 166:39]
  wire  _GEN_34711 = io_i_ex_res_packs_0_valid ? _GEN_32535 : _GEN_30293; // @[rob.scala 166:39]
  wire  _GEN_34712 = io_i_ex_res_packs_0_valid ? _GEN_32536 : _GEN_30294; // @[rob.scala 166:39]
  wire  _GEN_34713 = io_i_ex_res_packs_0_valid ? _GEN_32537 : _GEN_30295; // @[rob.scala 166:39]
  wire  _GEN_34714 = io_i_ex_res_packs_0_valid ? _GEN_32538 : _GEN_30296; // @[rob.scala 166:39]
  wire  _GEN_34715 = io_i_ex_res_packs_0_valid ? _GEN_32539 : _GEN_30297; // @[rob.scala 166:39]
  wire  _GEN_34716 = io_i_ex_res_packs_0_valid ? _GEN_32540 : _GEN_30298; // @[rob.scala 166:39]
  wire  _GEN_34717 = io_i_ex_res_packs_0_valid ? _GEN_32541 : _GEN_30299; // @[rob.scala 166:39]
  wire  _GEN_34718 = io_i_ex_res_packs_0_valid ? _GEN_32542 : _GEN_30300; // @[rob.scala 166:39]
  wire  _GEN_34719 = io_i_ex_res_packs_0_valid ? _GEN_32543 : _GEN_30301; // @[rob.scala 166:39]
  wire  _GEN_34720 = io_i_ex_res_packs_0_valid ? _GEN_32544 : _GEN_30302; // @[rob.scala 166:39]
  wire  _GEN_34721 = io_i_ex_res_packs_0_valid ? _GEN_32545 : _GEN_30303; // @[rob.scala 166:39]
  wire  _GEN_34722 = io_i_ex_res_packs_0_valid ? _GEN_32546 : _GEN_30304; // @[rob.scala 166:39]
  wire  _GEN_34723 = io_i_ex_res_packs_0_valid ? _GEN_32547 : _GEN_30305; // @[rob.scala 166:39]
  wire  _GEN_34724 = io_i_ex_res_packs_0_valid ? _GEN_32548 : _GEN_30306; // @[rob.scala 166:39]
  wire  _GEN_34725 = io_i_ex_res_packs_0_valid ? _GEN_32549 : _GEN_30307; // @[rob.scala 166:39]
  wire  _GEN_34726 = io_i_ex_res_packs_0_valid ? _GEN_32550 : _GEN_30308; // @[rob.scala 166:39]
  wire  _GEN_34727 = io_i_ex_res_packs_0_valid ? _GEN_32551 : _GEN_30309; // @[rob.scala 166:39]
  wire  _GEN_34728 = io_i_ex_res_packs_0_valid ? _GEN_32552 : _GEN_30310; // @[rob.scala 166:39]
  wire  _GEN_34729 = io_i_ex_res_packs_0_valid ? _GEN_32553 : _GEN_30311; // @[rob.scala 166:39]
  wire  _GEN_34730 = io_i_ex_res_packs_0_valid ? _GEN_32554 : _GEN_30312; // @[rob.scala 166:39]
  wire  _GEN_34731 = io_i_ex_res_packs_0_valid ? _GEN_32555 : _GEN_30313; // @[rob.scala 166:39]
  wire  _GEN_34732 = io_i_ex_res_packs_0_valid ? _GEN_32556 : _GEN_30314; // @[rob.scala 166:39]
  wire  _GEN_34733 = io_i_ex_res_packs_0_valid ? _GEN_32557 : _GEN_30315; // @[rob.scala 166:39]
  wire  _GEN_34734 = io_i_ex_res_packs_0_valid ? _GEN_32558 : _GEN_30316; // @[rob.scala 166:39]
  wire  _GEN_34735 = io_i_ex_res_packs_0_valid ? _GEN_32559 : _GEN_30317; // @[rob.scala 166:39]
  wire  _GEN_34736 = io_i_ex_res_packs_0_valid ? _GEN_32560 : _GEN_30318; // @[rob.scala 166:39]
  wire  _GEN_34737 = io_i_ex_res_packs_0_valid ? _GEN_32561 : _GEN_30319; // @[rob.scala 166:39]
  wire  _GEN_34738 = io_i_ex_res_packs_0_valid ? _GEN_32562 : _GEN_30320; // @[rob.scala 166:39]
  wire  _GEN_34739 = io_i_ex_res_packs_0_valid ? _GEN_32563 : _GEN_30321; // @[rob.scala 166:39]
  wire  _GEN_34740 = io_i_ex_res_packs_0_valid ? _GEN_32564 : _GEN_30322; // @[rob.scala 166:39]
  wire  _GEN_34741 = io_i_ex_res_packs_0_valid ? _GEN_32565 : _GEN_30323; // @[rob.scala 166:39]
  wire  _GEN_34742 = io_i_ex_res_packs_0_valid ? _GEN_32566 : _GEN_30324; // @[rob.scala 166:39]
  wire  _GEN_34743 = io_i_ex_res_packs_0_valid ? _GEN_32567 : _GEN_30325; // @[rob.scala 166:39]
  wire  _GEN_34744 = io_i_ex_res_packs_0_valid ? _GEN_32568 : _GEN_30326; // @[rob.scala 166:39]
  wire  _GEN_34745 = io_i_ex_res_packs_0_valid ? _GEN_32569 : _GEN_30327; // @[rob.scala 166:39]
  wire  _GEN_34746 = io_i_ex_res_packs_0_valid ? _GEN_32570 : _GEN_30328; // @[rob.scala 166:39]
  wire  _GEN_34747 = io_i_ex_res_packs_0_valid ? _GEN_32571 : _GEN_30329; // @[rob.scala 166:39]
  wire  _GEN_34748 = io_i_ex_res_packs_0_valid ? _GEN_32572 : _GEN_30330; // @[rob.scala 166:39]
  wire  _GEN_34749 = io_i_ex_res_packs_0_valid ? _GEN_32573 : _GEN_30331; // @[rob.scala 166:39]
  wire  _GEN_34750 = io_i_ex_res_packs_0_valid ? _GEN_32574 : _GEN_30332; // @[rob.scala 166:39]
  wire  _GEN_34751 = io_i_ex_res_packs_0_valid ? _GEN_32575 : _GEN_30333; // @[rob.scala 166:39]
  wire  _GEN_34752 = io_i_ex_res_packs_0_valid ? _GEN_32576 : _GEN_30334; // @[rob.scala 166:39]
  wire  _GEN_34753 = io_i_ex_res_packs_0_valid ? _GEN_32577 : _GEN_30335; // @[rob.scala 166:39]
  wire  _GEN_34754 = io_i_ex_res_packs_0_valid ? _GEN_32578 : _GEN_30336; // @[rob.scala 166:39]
  wire  _GEN_34755 = io_i_ex_res_packs_0_valid ? _GEN_32579 : _GEN_30337; // @[rob.scala 166:39]
  wire  _GEN_34756 = io_i_ex_res_packs_0_valid ? _GEN_32580 : _GEN_30338; // @[rob.scala 166:39]
  wire  _GEN_34757 = io_i_ex_res_packs_0_valid ? _GEN_32581 : _GEN_30339; // @[rob.scala 166:39]
  wire  _GEN_34758 = _GEN_42193 | _GEN_32582; // @[rob.scala 173:{53,53}]
  wire  _GEN_34759 = _GEN_42194 | _GEN_32583; // @[rob.scala 173:{53,53}]
  wire  _GEN_34760 = _GEN_42195 | _GEN_32584; // @[rob.scala 173:{53,53}]
  wire  _GEN_34761 = _GEN_42196 | _GEN_32585; // @[rob.scala 173:{53,53}]
  wire  _GEN_34762 = _GEN_42197 | _GEN_32586; // @[rob.scala 173:{53,53}]
  wire  _GEN_34763 = _GEN_42198 | _GEN_32587; // @[rob.scala 173:{53,53}]
  wire  _GEN_34764 = _GEN_42199 | _GEN_32588; // @[rob.scala 173:{53,53}]
  wire  _GEN_34765 = _GEN_42200 | _GEN_32589; // @[rob.scala 173:{53,53}]
  wire  _GEN_34766 = _GEN_42201 | _GEN_32590; // @[rob.scala 173:{53,53}]
  wire  _GEN_34767 = _GEN_42202 | _GEN_32591; // @[rob.scala 173:{53,53}]
  wire  _GEN_34768 = _GEN_42203 | _GEN_32592; // @[rob.scala 173:{53,53}]
  wire  _GEN_34769 = _GEN_42204 | _GEN_32593; // @[rob.scala 173:{53,53}]
  wire  _GEN_34770 = _GEN_42205 | _GEN_32594; // @[rob.scala 173:{53,53}]
  wire  _GEN_34771 = _GEN_42206 | _GEN_32595; // @[rob.scala 173:{53,53}]
  wire  _GEN_34772 = _GEN_42207 | _GEN_32596; // @[rob.scala 173:{53,53}]
  wire  _GEN_34773 = _GEN_42208 | _GEN_32597; // @[rob.scala 173:{53,53}]
  wire  _GEN_34774 = _GEN_42209 | _GEN_32598; // @[rob.scala 173:{53,53}]
  wire  _GEN_34775 = _GEN_42210 | _GEN_32599; // @[rob.scala 173:{53,53}]
  wire  _GEN_34776 = _GEN_42211 | _GEN_32600; // @[rob.scala 173:{53,53}]
  wire  _GEN_34777 = _GEN_42212 | _GEN_32601; // @[rob.scala 173:{53,53}]
  wire  _GEN_34778 = _GEN_42213 | _GEN_32602; // @[rob.scala 173:{53,53}]
  wire  _GEN_34779 = _GEN_42214 | _GEN_32603; // @[rob.scala 173:{53,53}]
  wire  _GEN_34780 = _GEN_42215 | _GEN_32604; // @[rob.scala 173:{53,53}]
  wire  _GEN_34781 = _GEN_42216 | _GEN_32605; // @[rob.scala 173:{53,53}]
  wire  _GEN_34782 = _GEN_42217 | _GEN_32606; // @[rob.scala 173:{53,53}]
  wire  _GEN_34783 = _GEN_42218 | _GEN_32607; // @[rob.scala 173:{53,53}]
  wire  _GEN_34784 = _GEN_42219 | _GEN_32608; // @[rob.scala 173:{53,53}]
  wire  _GEN_34785 = _GEN_42220 | _GEN_32609; // @[rob.scala 173:{53,53}]
  wire  _GEN_34786 = _GEN_42221 | _GEN_32610; // @[rob.scala 173:{53,53}]
  wire  _GEN_34787 = _GEN_42222 | _GEN_32611; // @[rob.scala 173:{53,53}]
  wire  _GEN_34788 = _GEN_42223 | _GEN_32612; // @[rob.scala 173:{53,53}]
  wire  _GEN_34789 = _GEN_42224 | _GEN_32613; // @[rob.scala 173:{53,53}]
  wire  _GEN_34790 = _GEN_42225 | _GEN_32614; // @[rob.scala 173:{53,53}]
  wire  _GEN_34791 = _GEN_42226 | _GEN_32615; // @[rob.scala 173:{53,53}]
  wire  _GEN_34792 = _GEN_42227 | _GEN_32616; // @[rob.scala 173:{53,53}]
  wire  _GEN_34793 = _GEN_42228 | _GEN_32617; // @[rob.scala 173:{53,53}]
  wire  _GEN_34794 = _GEN_42229 | _GEN_32618; // @[rob.scala 173:{53,53}]
  wire  _GEN_34795 = _GEN_42230 | _GEN_32619; // @[rob.scala 173:{53,53}]
  wire  _GEN_34796 = _GEN_42231 | _GEN_32620; // @[rob.scala 173:{53,53}]
  wire  _GEN_34797 = _GEN_42232 | _GEN_32621; // @[rob.scala 173:{53,53}]
  wire  _GEN_34798 = _GEN_42233 | _GEN_32622; // @[rob.scala 173:{53,53}]
  wire  _GEN_34799 = _GEN_42234 | _GEN_32623; // @[rob.scala 173:{53,53}]
  wire  _GEN_34800 = _GEN_42235 | _GEN_32624; // @[rob.scala 173:{53,53}]
  wire  _GEN_34801 = _GEN_42236 | _GEN_32625; // @[rob.scala 173:{53,53}]
  wire  _GEN_34802 = _GEN_42237 | _GEN_32626; // @[rob.scala 173:{53,53}]
  wire  _GEN_34803 = _GEN_42238 | _GEN_32627; // @[rob.scala 173:{53,53}]
  wire  _GEN_34804 = _GEN_42239 | _GEN_32628; // @[rob.scala 173:{53,53}]
  wire  _GEN_34805 = _GEN_42240 | _GEN_32629; // @[rob.scala 173:{53,53}]
  wire  _GEN_34806 = _GEN_42241 | _GEN_32630; // @[rob.scala 173:{53,53}]
  wire  _GEN_34807 = _GEN_42242 | _GEN_32631; // @[rob.scala 173:{53,53}]
  wire  _GEN_34808 = _GEN_42243 | _GEN_32632; // @[rob.scala 173:{53,53}]
  wire  _GEN_34809 = _GEN_42244 | _GEN_32633; // @[rob.scala 173:{53,53}]
  wire  _GEN_34810 = _GEN_42245 | _GEN_32634; // @[rob.scala 173:{53,53}]
  wire  _GEN_34811 = _GEN_42246 | _GEN_32635; // @[rob.scala 173:{53,53}]
  wire  _GEN_34812 = _GEN_42247 | _GEN_32636; // @[rob.scala 173:{53,53}]
  wire  _GEN_34813 = _GEN_42248 | _GEN_32637; // @[rob.scala 173:{53,53}]
  wire  _GEN_34814 = _GEN_42249 | _GEN_32638; // @[rob.scala 173:{53,53}]
  wire  _GEN_34815 = _GEN_42250 | _GEN_32639; // @[rob.scala 173:{53,53}]
  wire  _GEN_34816 = _GEN_42251 | _GEN_32640; // @[rob.scala 173:{53,53}]
  wire  _GEN_34817 = _GEN_42252 | _GEN_32641; // @[rob.scala 173:{53,53}]
  wire  _GEN_34818 = _GEN_42253 | _GEN_32642; // @[rob.scala 173:{53,53}]
  wire  _GEN_34819 = _GEN_42254 | _GEN_32643; // @[rob.scala 173:{53,53}]
  wire  _GEN_34820 = _GEN_42255 | _GEN_32644; // @[rob.scala 173:{53,53}]
  wire  _GEN_34821 = _GEN_42256 | _GEN_32645; // @[rob.scala 173:{53,53}]
  wire  _GEN_36870 = _GEN_42193 | _GEN_34694; // @[rob.scala 176:{52,52}]
  wire  _GEN_36871 = _GEN_42194 | _GEN_34695; // @[rob.scala 176:{52,52}]
  wire  _GEN_36872 = _GEN_42195 | _GEN_34696; // @[rob.scala 176:{52,52}]
  wire  _GEN_36873 = _GEN_42196 | _GEN_34697; // @[rob.scala 176:{52,52}]
  wire  _GEN_36874 = _GEN_42197 | _GEN_34698; // @[rob.scala 176:{52,52}]
  wire  _GEN_36875 = _GEN_42198 | _GEN_34699; // @[rob.scala 176:{52,52}]
  wire  _GEN_36876 = _GEN_42199 | _GEN_34700; // @[rob.scala 176:{52,52}]
  wire  _GEN_36877 = _GEN_42200 | _GEN_34701; // @[rob.scala 176:{52,52}]
  wire  _GEN_36878 = _GEN_42201 | _GEN_34702; // @[rob.scala 176:{52,52}]
  wire  _GEN_36879 = _GEN_42202 | _GEN_34703; // @[rob.scala 176:{52,52}]
  wire  _GEN_36880 = _GEN_42203 | _GEN_34704; // @[rob.scala 176:{52,52}]
  wire  _GEN_36881 = _GEN_42204 | _GEN_34705; // @[rob.scala 176:{52,52}]
  wire  _GEN_36882 = _GEN_42205 | _GEN_34706; // @[rob.scala 176:{52,52}]
  wire  _GEN_36883 = _GEN_42206 | _GEN_34707; // @[rob.scala 176:{52,52}]
  wire  _GEN_36884 = _GEN_42207 | _GEN_34708; // @[rob.scala 176:{52,52}]
  wire  _GEN_36885 = _GEN_42208 | _GEN_34709; // @[rob.scala 176:{52,52}]
  wire  _GEN_36886 = _GEN_42209 | _GEN_34710; // @[rob.scala 176:{52,52}]
  wire  _GEN_36887 = _GEN_42210 | _GEN_34711; // @[rob.scala 176:{52,52}]
  wire  _GEN_36888 = _GEN_42211 | _GEN_34712; // @[rob.scala 176:{52,52}]
  wire  _GEN_36889 = _GEN_42212 | _GEN_34713; // @[rob.scala 176:{52,52}]
  wire  _GEN_36890 = _GEN_42213 | _GEN_34714; // @[rob.scala 176:{52,52}]
  wire  _GEN_36891 = _GEN_42214 | _GEN_34715; // @[rob.scala 176:{52,52}]
  wire  _GEN_36892 = _GEN_42215 | _GEN_34716; // @[rob.scala 176:{52,52}]
  wire  _GEN_36893 = _GEN_42216 | _GEN_34717; // @[rob.scala 176:{52,52}]
  wire  _GEN_36894 = _GEN_42217 | _GEN_34718; // @[rob.scala 176:{52,52}]
  wire  _GEN_36895 = _GEN_42218 | _GEN_34719; // @[rob.scala 176:{52,52}]
  wire  _GEN_36896 = _GEN_42219 | _GEN_34720; // @[rob.scala 176:{52,52}]
  wire  _GEN_36897 = _GEN_42220 | _GEN_34721; // @[rob.scala 176:{52,52}]
  wire  _GEN_36898 = _GEN_42221 | _GEN_34722; // @[rob.scala 176:{52,52}]
  wire  _GEN_36899 = _GEN_42222 | _GEN_34723; // @[rob.scala 176:{52,52}]
  wire  _GEN_36900 = _GEN_42223 | _GEN_34724; // @[rob.scala 176:{52,52}]
  wire  _GEN_36901 = _GEN_42224 | _GEN_34725; // @[rob.scala 176:{52,52}]
  wire  _GEN_36902 = _GEN_42225 | _GEN_34726; // @[rob.scala 176:{52,52}]
  wire  _GEN_36903 = _GEN_42226 | _GEN_34727; // @[rob.scala 176:{52,52}]
  wire  _GEN_36904 = _GEN_42227 | _GEN_34728; // @[rob.scala 176:{52,52}]
  wire  _GEN_36905 = _GEN_42228 | _GEN_34729; // @[rob.scala 176:{52,52}]
  wire  _GEN_36906 = _GEN_42229 | _GEN_34730; // @[rob.scala 176:{52,52}]
  wire  _GEN_36907 = _GEN_42230 | _GEN_34731; // @[rob.scala 176:{52,52}]
  wire  _GEN_36908 = _GEN_42231 | _GEN_34732; // @[rob.scala 176:{52,52}]
  wire  _GEN_36909 = _GEN_42232 | _GEN_34733; // @[rob.scala 176:{52,52}]
  wire  _GEN_36910 = _GEN_42233 | _GEN_34734; // @[rob.scala 176:{52,52}]
  wire  _GEN_36911 = _GEN_42234 | _GEN_34735; // @[rob.scala 176:{52,52}]
  wire  _GEN_36912 = _GEN_42235 | _GEN_34736; // @[rob.scala 176:{52,52}]
  wire  _GEN_36913 = _GEN_42236 | _GEN_34737; // @[rob.scala 176:{52,52}]
  wire  _GEN_36914 = _GEN_42237 | _GEN_34738; // @[rob.scala 176:{52,52}]
  wire  _GEN_36915 = _GEN_42238 | _GEN_34739; // @[rob.scala 176:{52,52}]
  wire  _GEN_36916 = _GEN_42239 | _GEN_34740; // @[rob.scala 176:{52,52}]
  wire  _GEN_36917 = _GEN_42240 | _GEN_34741; // @[rob.scala 176:{52,52}]
  wire  _GEN_36918 = _GEN_42241 | _GEN_34742; // @[rob.scala 176:{52,52}]
  wire  _GEN_36919 = _GEN_42242 | _GEN_34743; // @[rob.scala 176:{52,52}]
  wire  _GEN_36920 = _GEN_42243 | _GEN_34744; // @[rob.scala 176:{52,52}]
  wire  _GEN_36921 = _GEN_42244 | _GEN_34745; // @[rob.scala 176:{52,52}]
  wire  _GEN_36922 = _GEN_42245 | _GEN_34746; // @[rob.scala 176:{52,52}]
  wire  _GEN_36923 = _GEN_42246 | _GEN_34747; // @[rob.scala 176:{52,52}]
  wire  _GEN_36924 = _GEN_42247 | _GEN_34748; // @[rob.scala 176:{52,52}]
  wire  _GEN_36925 = _GEN_42248 | _GEN_34749; // @[rob.scala 176:{52,52}]
  wire  _GEN_36926 = _GEN_42249 | _GEN_34750; // @[rob.scala 176:{52,52}]
  wire  _GEN_36927 = _GEN_42250 | _GEN_34751; // @[rob.scala 176:{52,52}]
  wire  _GEN_36928 = _GEN_42251 | _GEN_34752; // @[rob.scala 176:{52,52}]
  wire  _GEN_36929 = _GEN_42252 | _GEN_34753; // @[rob.scala 176:{52,52}]
  wire  _GEN_36930 = _GEN_42253 | _GEN_34754; // @[rob.scala 176:{52,52}]
  wire  _GEN_36931 = _GEN_42254 | _GEN_34755; // @[rob.scala 176:{52,52}]
  wire  _GEN_36932 = _GEN_42255 | _GEN_34756; // @[rob.scala 176:{52,52}]
  wire  _GEN_36933 = _GEN_42256 | _GEN_34757; // @[rob.scala 176:{52,52}]
  wire  _GEN_36934 = io_i_ex_res_packs_1_valid ? _GEN_34758 : _GEN_32582; // @[rob.scala 172:39]
  wire  _GEN_36935 = io_i_ex_res_packs_1_valid ? _GEN_34759 : _GEN_32583; // @[rob.scala 172:39]
  wire  _GEN_36936 = io_i_ex_res_packs_1_valid ? _GEN_34760 : _GEN_32584; // @[rob.scala 172:39]
  wire  _GEN_36937 = io_i_ex_res_packs_1_valid ? _GEN_34761 : _GEN_32585; // @[rob.scala 172:39]
  wire  _GEN_36938 = io_i_ex_res_packs_1_valid ? _GEN_34762 : _GEN_32586; // @[rob.scala 172:39]
  wire  _GEN_36939 = io_i_ex_res_packs_1_valid ? _GEN_34763 : _GEN_32587; // @[rob.scala 172:39]
  wire  _GEN_36940 = io_i_ex_res_packs_1_valid ? _GEN_34764 : _GEN_32588; // @[rob.scala 172:39]
  wire  _GEN_36941 = io_i_ex_res_packs_1_valid ? _GEN_34765 : _GEN_32589; // @[rob.scala 172:39]
  wire  _GEN_36942 = io_i_ex_res_packs_1_valid ? _GEN_34766 : _GEN_32590; // @[rob.scala 172:39]
  wire  _GEN_36943 = io_i_ex_res_packs_1_valid ? _GEN_34767 : _GEN_32591; // @[rob.scala 172:39]
  wire  _GEN_36944 = io_i_ex_res_packs_1_valid ? _GEN_34768 : _GEN_32592; // @[rob.scala 172:39]
  wire  _GEN_36945 = io_i_ex_res_packs_1_valid ? _GEN_34769 : _GEN_32593; // @[rob.scala 172:39]
  wire  _GEN_36946 = io_i_ex_res_packs_1_valid ? _GEN_34770 : _GEN_32594; // @[rob.scala 172:39]
  wire  _GEN_36947 = io_i_ex_res_packs_1_valid ? _GEN_34771 : _GEN_32595; // @[rob.scala 172:39]
  wire  _GEN_36948 = io_i_ex_res_packs_1_valid ? _GEN_34772 : _GEN_32596; // @[rob.scala 172:39]
  wire  _GEN_36949 = io_i_ex_res_packs_1_valid ? _GEN_34773 : _GEN_32597; // @[rob.scala 172:39]
  wire  _GEN_36950 = io_i_ex_res_packs_1_valid ? _GEN_34774 : _GEN_32598; // @[rob.scala 172:39]
  wire  _GEN_36951 = io_i_ex_res_packs_1_valid ? _GEN_34775 : _GEN_32599; // @[rob.scala 172:39]
  wire  _GEN_36952 = io_i_ex_res_packs_1_valid ? _GEN_34776 : _GEN_32600; // @[rob.scala 172:39]
  wire  _GEN_36953 = io_i_ex_res_packs_1_valid ? _GEN_34777 : _GEN_32601; // @[rob.scala 172:39]
  wire  _GEN_36954 = io_i_ex_res_packs_1_valid ? _GEN_34778 : _GEN_32602; // @[rob.scala 172:39]
  wire  _GEN_36955 = io_i_ex_res_packs_1_valid ? _GEN_34779 : _GEN_32603; // @[rob.scala 172:39]
  wire  _GEN_36956 = io_i_ex_res_packs_1_valid ? _GEN_34780 : _GEN_32604; // @[rob.scala 172:39]
  wire  _GEN_36957 = io_i_ex_res_packs_1_valid ? _GEN_34781 : _GEN_32605; // @[rob.scala 172:39]
  wire  _GEN_36958 = io_i_ex_res_packs_1_valid ? _GEN_34782 : _GEN_32606; // @[rob.scala 172:39]
  wire  _GEN_36959 = io_i_ex_res_packs_1_valid ? _GEN_34783 : _GEN_32607; // @[rob.scala 172:39]
  wire  _GEN_36960 = io_i_ex_res_packs_1_valid ? _GEN_34784 : _GEN_32608; // @[rob.scala 172:39]
  wire  _GEN_36961 = io_i_ex_res_packs_1_valid ? _GEN_34785 : _GEN_32609; // @[rob.scala 172:39]
  wire  _GEN_36962 = io_i_ex_res_packs_1_valid ? _GEN_34786 : _GEN_32610; // @[rob.scala 172:39]
  wire  _GEN_36963 = io_i_ex_res_packs_1_valid ? _GEN_34787 : _GEN_32611; // @[rob.scala 172:39]
  wire  _GEN_36964 = io_i_ex_res_packs_1_valid ? _GEN_34788 : _GEN_32612; // @[rob.scala 172:39]
  wire  _GEN_36965 = io_i_ex_res_packs_1_valid ? _GEN_34789 : _GEN_32613; // @[rob.scala 172:39]
  wire  _GEN_36966 = io_i_ex_res_packs_1_valid ? _GEN_34790 : _GEN_32614; // @[rob.scala 172:39]
  wire  _GEN_36967 = io_i_ex_res_packs_1_valid ? _GEN_34791 : _GEN_32615; // @[rob.scala 172:39]
  wire  _GEN_36968 = io_i_ex_res_packs_1_valid ? _GEN_34792 : _GEN_32616; // @[rob.scala 172:39]
  wire  _GEN_36969 = io_i_ex_res_packs_1_valid ? _GEN_34793 : _GEN_32617; // @[rob.scala 172:39]
  wire  _GEN_36970 = io_i_ex_res_packs_1_valid ? _GEN_34794 : _GEN_32618; // @[rob.scala 172:39]
  wire  _GEN_36971 = io_i_ex_res_packs_1_valid ? _GEN_34795 : _GEN_32619; // @[rob.scala 172:39]
  wire  _GEN_36972 = io_i_ex_res_packs_1_valid ? _GEN_34796 : _GEN_32620; // @[rob.scala 172:39]
  wire  _GEN_36973 = io_i_ex_res_packs_1_valid ? _GEN_34797 : _GEN_32621; // @[rob.scala 172:39]
  wire  _GEN_36974 = io_i_ex_res_packs_1_valid ? _GEN_34798 : _GEN_32622; // @[rob.scala 172:39]
  wire  _GEN_36975 = io_i_ex_res_packs_1_valid ? _GEN_34799 : _GEN_32623; // @[rob.scala 172:39]
  wire  _GEN_36976 = io_i_ex_res_packs_1_valid ? _GEN_34800 : _GEN_32624; // @[rob.scala 172:39]
  wire  _GEN_36977 = io_i_ex_res_packs_1_valid ? _GEN_34801 : _GEN_32625; // @[rob.scala 172:39]
  wire  _GEN_36978 = io_i_ex_res_packs_1_valid ? _GEN_34802 : _GEN_32626; // @[rob.scala 172:39]
  wire  _GEN_36979 = io_i_ex_res_packs_1_valid ? _GEN_34803 : _GEN_32627; // @[rob.scala 172:39]
  wire  _GEN_36980 = io_i_ex_res_packs_1_valid ? _GEN_34804 : _GEN_32628; // @[rob.scala 172:39]
  wire  _GEN_36981 = io_i_ex_res_packs_1_valid ? _GEN_34805 : _GEN_32629; // @[rob.scala 172:39]
  wire  _GEN_36982 = io_i_ex_res_packs_1_valid ? _GEN_34806 : _GEN_32630; // @[rob.scala 172:39]
  wire  _GEN_36983 = io_i_ex_res_packs_1_valid ? _GEN_34807 : _GEN_32631; // @[rob.scala 172:39]
  wire  _GEN_36984 = io_i_ex_res_packs_1_valid ? _GEN_34808 : _GEN_32632; // @[rob.scala 172:39]
  wire  _GEN_36985 = io_i_ex_res_packs_1_valid ? _GEN_34809 : _GEN_32633; // @[rob.scala 172:39]
  wire  _GEN_36986 = io_i_ex_res_packs_1_valid ? _GEN_34810 : _GEN_32634; // @[rob.scala 172:39]
  wire  _GEN_36987 = io_i_ex_res_packs_1_valid ? _GEN_34811 : _GEN_32635; // @[rob.scala 172:39]
  wire  _GEN_36988 = io_i_ex_res_packs_1_valid ? _GEN_34812 : _GEN_32636; // @[rob.scala 172:39]
  wire  _GEN_36989 = io_i_ex_res_packs_1_valid ? _GEN_34813 : _GEN_32637; // @[rob.scala 172:39]
  wire  _GEN_36990 = io_i_ex_res_packs_1_valid ? _GEN_34814 : _GEN_32638; // @[rob.scala 172:39]
  wire  _GEN_36991 = io_i_ex_res_packs_1_valid ? _GEN_34815 : _GEN_32639; // @[rob.scala 172:39]
  wire  _GEN_36992 = io_i_ex_res_packs_1_valid ? _GEN_34816 : _GEN_32640; // @[rob.scala 172:39]
  wire  _GEN_36993 = io_i_ex_res_packs_1_valid ? _GEN_34817 : _GEN_32641; // @[rob.scala 172:39]
  wire  _GEN_36994 = io_i_ex_res_packs_1_valid ? _GEN_34818 : _GEN_32642; // @[rob.scala 172:39]
  wire  _GEN_36995 = io_i_ex_res_packs_1_valid ? _GEN_34819 : _GEN_32643; // @[rob.scala 172:39]
  wire  _GEN_36996 = io_i_ex_res_packs_1_valid ? _GEN_34820 : _GEN_32644; // @[rob.scala 172:39]
  wire  _GEN_36997 = io_i_ex_res_packs_1_valid ? _GEN_34821 : _GEN_32645; // @[rob.scala 172:39]
  wire  _GEN_39110 = 6'h0 == commit_ptr[5:0] ? 1'h0 : _GEN_36934; // @[rob.scala 180:{31,31}]
  wire  _GEN_39111 = 6'h1 == commit_ptr[5:0] ? 1'h0 : _GEN_36935; // @[rob.scala 180:{31,31}]
  wire  _GEN_39112 = 6'h2 == commit_ptr[5:0] ? 1'h0 : _GEN_36936; // @[rob.scala 180:{31,31}]
  wire  _GEN_39113 = 6'h3 == commit_ptr[5:0] ? 1'h0 : _GEN_36937; // @[rob.scala 180:{31,31}]
  wire  _GEN_39114 = 6'h4 == commit_ptr[5:0] ? 1'h0 : _GEN_36938; // @[rob.scala 180:{31,31}]
  wire  _GEN_39115 = 6'h5 == commit_ptr[5:0] ? 1'h0 : _GEN_36939; // @[rob.scala 180:{31,31}]
  wire  _GEN_39116 = 6'h6 == commit_ptr[5:0] ? 1'h0 : _GEN_36940; // @[rob.scala 180:{31,31}]
  wire  _GEN_39117 = 6'h7 == commit_ptr[5:0] ? 1'h0 : _GEN_36941; // @[rob.scala 180:{31,31}]
  wire  _GEN_39118 = 6'h8 == commit_ptr[5:0] ? 1'h0 : _GEN_36942; // @[rob.scala 180:{31,31}]
  wire  _GEN_39119 = 6'h9 == commit_ptr[5:0] ? 1'h0 : _GEN_36943; // @[rob.scala 180:{31,31}]
  wire  _GEN_39120 = 6'ha == commit_ptr[5:0] ? 1'h0 : _GEN_36944; // @[rob.scala 180:{31,31}]
  wire  _GEN_39121 = 6'hb == commit_ptr[5:0] ? 1'h0 : _GEN_36945; // @[rob.scala 180:{31,31}]
  wire  _GEN_39122 = 6'hc == commit_ptr[5:0] ? 1'h0 : _GEN_36946; // @[rob.scala 180:{31,31}]
  wire  _GEN_39123 = 6'hd == commit_ptr[5:0] ? 1'h0 : _GEN_36947; // @[rob.scala 180:{31,31}]
  wire  _GEN_39124 = 6'he == commit_ptr[5:0] ? 1'h0 : _GEN_36948; // @[rob.scala 180:{31,31}]
  wire  _GEN_39125 = 6'hf == commit_ptr[5:0] ? 1'h0 : _GEN_36949; // @[rob.scala 180:{31,31}]
  wire  _GEN_39126 = 6'h10 == commit_ptr[5:0] ? 1'h0 : _GEN_36950; // @[rob.scala 180:{31,31}]
  wire  _GEN_39127 = 6'h11 == commit_ptr[5:0] ? 1'h0 : _GEN_36951; // @[rob.scala 180:{31,31}]
  wire  _GEN_39128 = 6'h12 == commit_ptr[5:0] ? 1'h0 : _GEN_36952; // @[rob.scala 180:{31,31}]
  wire  _GEN_39129 = 6'h13 == commit_ptr[5:0] ? 1'h0 : _GEN_36953; // @[rob.scala 180:{31,31}]
  wire  _GEN_39130 = 6'h14 == commit_ptr[5:0] ? 1'h0 : _GEN_36954; // @[rob.scala 180:{31,31}]
  wire  _GEN_39131 = 6'h15 == commit_ptr[5:0] ? 1'h0 : _GEN_36955; // @[rob.scala 180:{31,31}]
  wire  _GEN_39132 = 6'h16 == commit_ptr[5:0] ? 1'h0 : _GEN_36956; // @[rob.scala 180:{31,31}]
  wire  _GEN_39133 = 6'h17 == commit_ptr[5:0] ? 1'h0 : _GEN_36957; // @[rob.scala 180:{31,31}]
  wire  _GEN_39134 = 6'h18 == commit_ptr[5:0] ? 1'h0 : _GEN_36958; // @[rob.scala 180:{31,31}]
  wire  _GEN_39135 = 6'h19 == commit_ptr[5:0] ? 1'h0 : _GEN_36959; // @[rob.scala 180:{31,31}]
  wire  _GEN_39136 = 6'h1a == commit_ptr[5:0] ? 1'h0 : _GEN_36960; // @[rob.scala 180:{31,31}]
  wire  _GEN_39137 = 6'h1b == commit_ptr[5:0] ? 1'h0 : _GEN_36961; // @[rob.scala 180:{31,31}]
  wire  _GEN_39138 = 6'h1c == commit_ptr[5:0] ? 1'h0 : _GEN_36962; // @[rob.scala 180:{31,31}]
  wire  _GEN_39139 = 6'h1d == commit_ptr[5:0] ? 1'h0 : _GEN_36963; // @[rob.scala 180:{31,31}]
  wire  _GEN_39140 = 6'h1e == commit_ptr[5:0] ? 1'h0 : _GEN_36964; // @[rob.scala 180:{31,31}]
  wire  _GEN_39141 = 6'h1f == commit_ptr[5:0] ? 1'h0 : _GEN_36965; // @[rob.scala 180:{31,31}]
  wire  _GEN_39142 = 6'h20 == commit_ptr[5:0] ? 1'h0 : _GEN_36966; // @[rob.scala 180:{31,31}]
  wire  _GEN_39143 = 6'h21 == commit_ptr[5:0] ? 1'h0 : _GEN_36967; // @[rob.scala 180:{31,31}]
  wire  _GEN_39144 = 6'h22 == commit_ptr[5:0] ? 1'h0 : _GEN_36968; // @[rob.scala 180:{31,31}]
  wire  _GEN_39145 = 6'h23 == commit_ptr[5:0] ? 1'h0 : _GEN_36969; // @[rob.scala 180:{31,31}]
  wire  _GEN_39146 = 6'h24 == commit_ptr[5:0] ? 1'h0 : _GEN_36970; // @[rob.scala 180:{31,31}]
  wire  _GEN_39147 = 6'h25 == commit_ptr[5:0] ? 1'h0 : _GEN_36971; // @[rob.scala 180:{31,31}]
  wire  _GEN_39148 = 6'h26 == commit_ptr[5:0] ? 1'h0 : _GEN_36972; // @[rob.scala 180:{31,31}]
  wire  _GEN_39149 = 6'h27 == commit_ptr[5:0] ? 1'h0 : _GEN_36973; // @[rob.scala 180:{31,31}]
  wire  _GEN_39150 = 6'h28 == commit_ptr[5:0] ? 1'h0 : _GEN_36974; // @[rob.scala 180:{31,31}]
  wire  _GEN_39151 = 6'h29 == commit_ptr[5:0] ? 1'h0 : _GEN_36975; // @[rob.scala 180:{31,31}]
  wire  _GEN_39152 = 6'h2a == commit_ptr[5:0] ? 1'h0 : _GEN_36976; // @[rob.scala 180:{31,31}]
  wire  _GEN_39153 = 6'h2b == commit_ptr[5:0] ? 1'h0 : _GEN_36977; // @[rob.scala 180:{31,31}]
  wire  _GEN_39154 = 6'h2c == commit_ptr[5:0] ? 1'h0 : _GEN_36978; // @[rob.scala 180:{31,31}]
  wire  _GEN_39155 = 6'h2d == commit_ptr[5:0] ? 1'h0 : _GEN_36979; // @[rob.scala 180:{31,31}]
  wire  _GEN_39156 = 6'h2e == commit_ptr[5:0] ? 1'h0 : _GEN_36980; // @[rob.scala 180:{31,31}]
  wire  _GEN_39157 = 6'h2f == commit_ptr[5:0] ? 1'h0 : _GEN_36981; // @[rob.scala 180:{31,31}]
  wire  _GEN_39158 = 6'h30 == commit_ptr[5:0] ? 1'h0 : _GEN_36982; // @[rob.scala 180:{31,31}]
  wire  _GEN_39159 = 6'h31 == commit_ptr[5:0] ? 1'h0 : _GEN_36983; // @[rob.scala 180:{31,31}]
  wire  _GEN_39160 = 6'h32 == commit_ptr[5:0] ? 1'h0 : _GEN_36984; // @[rob.scala 180:{31,31}]
  wire  _GEN_39161 = 6'h33 == commit_ptr[5:0] ? 1'h0 : _GEN_36985; // @[rob.scala 180:{31,31}]
  wire  _GEN_39162 = 6'h34 == commit_ptr[5:0] ? 1'h0 : _GEN_36986; // @[rob.scala 180:{31,31}]
  wire  _GEN_39163 = 6'h35 == commit_ptr[5:0] ? 1'h0 : _GEN_36987; // @[rob.scala 180:{31,31}]
  wire  _GEN_39164 = 6'h36 == commit_ptr[5:0] ? 1'h0 : _GEN_36988; // @[rob.scala 180:{31,31}]
  wire  _GEN_39165 = 6'h37 == commit_ptr[5:0] ? 1'h0 : _GEN_36989; // @[rob.scala 180:{31,31}]
  wire  _GEN_39166 = 6'h38 == commit_ptr[5:0] ? 1'h0 : _GEN_36990; // @[rob.scala 180:{31,31}]
  wire  _GEN_39167 = 6'h39 == commit_ptr[5:0] ? 1'h0 : _GEN_36991; // @[rob.scala 180:{31,31}]
  wire  _GEN_39168 = 6'h3a == commit_ptr[5:0] ? 1'h0 : _GEN_36992; // @[rob.scala 180:{31,31}]
  wire  _GEN_39169 = 6'h3b == commit_ptr[5:0] ? 1'h0 : _GEN_36993; // @[rob.scala 180:{31,31}]
  wire  _GEN_39170 = 6'h3c == commit_ptr[5:0] ? 1'h0 : _GEN_36994; // @[rob.scala 180:{31,31}]
  wire  _GEN_39171 = 6'h3d == commit_ptr[5:0] ? 1'h0 : _GEN_36995; // @[rob.scala 180:{31,31}]
  wire  _GEN_39172 = 6'h3e == commit_ptr[5:0] ? 1'h0 : _GEN_36996; // @[rob.scala 180:{31,31}]
  wire  _GEN_39173 = 6'h3f == commit_ptr[5:0] ? 1'h0 : _GEN_36997; // @[rob.scala 180:{31,31}]
  wire  _GEN_39174 = 6'h0 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39110; // @[rob.scala 181:{35,35}]
  wire  _GEN_39175 = 6'h1 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39111; // @[rob.scala 181:{35,35}]
  wire  _GEN_39176 = 6'h2 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39112; // @[rob.scala 181:{35,35}]
  wire  _GEN_39177 = 6'h3 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39113; // @[rob.scala 181:{35,35}]
  wire  _GEN_39178 = 6'h4 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39114; // @[rob.scala 181:{35,35}]
  wire  _GEN_39179 = 6'h5 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39115; // @[rob.scala 181:{35,35}]
  wire  _GEN_39180 = 6'h6 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39116; // @[rob.scala 181:{35,35}]
  wire  _GEN_39181 = 6'h7 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39117; // @[rob.scala 181:{35,35}]
  wire  _GEN_39182 = 6'h8 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39118; // @[rob.scala 181:{35,35}]
  wire  _GEN_39183 = 6'h9 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39119; // @[rob.scala 181:{35,35}]
  wire  _GEN_39184 = 6'ha == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39120; // @[rob.scala 181:{35,35}]
  wire  _GEN_39185 = 6'hb == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39121; // @[rob.scala 181:{35,35}]
  wire  _GEN_39186 = 6'hc == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39122; // @[rob.scala 181:{35,35}]
  wire  _GEN_39187 = 6'hd == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39123; // @[rob.scala 181:{35,35}]
  wire  _GEN_39188 = 6'he == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39124; // @[rob.scala 181:{35,35}]
  wire  _GEN_39189 = 6'hf == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39125; // @[rob.scala 181:{35,35}]
  wire  _GEN_39190 = 6'h10 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39126; // @[rob.scala 181:{35,35}]
  wire  _GEN_39191 = 6'h11 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39127; // @[rob.scala 181:{35,35}]
  wire  _GEN_39192 = 6'h12 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39128; // @[rob.scala 181:{35,35}]
  wire  _GEN_39193 = 6'h13 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39129; // @[rob.scala 181:{35,35}]
  wire  _GEN_39194 = 6'h14 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39130; // @[rob.scala 181:{35,35}]
  wire  _GEN_39195 = 6'h15 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39131; // @[rob.scala 181:{35,35}]
  wire  _GEN_39196 = 6'h16 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39132; // @[rob.scala 181:{35,35}]
  wire  _GEN_39197 = 6'h17 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39133; // @[rob.scala 181:{35,35}]
  wire  _GEN_39198 = 6'h18 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39134; // @[rob.scala 181:{35,35}]
  wire  _GEN_39199 = 6'h19 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39135; // @[rob.scala 181:{35,35}]
  wire  _GEN_39200 = 6'h1a == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39136; // @[rob.scala 181:{35,35}]
  wire  _GEN_39201 = 6'h1b == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39137; // @[rob.scala 181:{35,35}]
  wire  _GEN_39202 = 6'h1c == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39138; // @[rob.scala 181:{35,35}]
  wire  _GEN_39203 = 6'h1d == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39139; // @[rob.scala 181:{35,35}]
  wire  _GEN_39204 = 6'h1e == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39140; // @[rob.scala 181:{35,35}]
  wire  _GEN_39205 = 6'h1f == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39141; // @[rob.scala 181:{35,35}]
  wire  _GEN_39206 = 6'h20 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39142; // @[rob.scala 181:{35,35}]
  wire  _GEN_39207 = 6'h21 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39143; // @[rob.scala 181:{35,35}]
  wire  _GEN_39208 = 6'h22 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39144; // @[rob.scala 181:{35,35}]
  wire  _GEN_39209 = 6'h23 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39145; // @[rob.scala 181:{35,35}]
  wire  _GEN_39210 = 6'h24 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39146; // @[rob.scala 181:{35,35}]
  wire  _GEN_39211 = 6'h25 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39147; // @[rob.scala 181:{35,35}]
  wire  _GEN_39212 = 6'h26 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39148; // @[rob.scala 181:{35,35}]
  wire  _GEN_39213 = 6'h27 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39149; // @[rob.scala 181:{35,35}]
  wire  _GEN_39214 = 6'h28 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39150; // @[rob.scala 181:{35,35}]
  wire  _GEN_39215 = 6'h29 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39151; // @[rob.scala 181:{35,35}]
  wire  _GEN_39216 = 6'h2a == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39152; // @[rob.scala 181:{35,35}]
  wire  _GEN_39217 = 6'h2b == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39153; // @[rob.scala 181:{35,35}]
  wire  _GEN_39218 = 6'h2c == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39154; // @[rob.scala 181:{35,35}]
  wire  _GEN_39219 = 6'h2d == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39155; // @[rob.scala 181:{35,35}]
  wire  _GEN_39220 = 6'h2e == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39156; // @[rob.scala 181:{35,35}]
  wire  _GEN_39221 = 6'h2f == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39157; // @[rob.scala 181:{35,35}]
  wire  _GEN_39222 = 6'h30 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39158; // @[rob.scala 181:{35,35}]
  wire  _GEN_39223 = 6'h31 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39159; // @[rob.scala 181:{35,35}]
  wire  _GEN_39224 = 6'h32 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39160; // @[rob.scala 181:{35,35}]
  wire  _GEN_39225 = 6'h33 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39161; // @[rob.scala 181:{35,35}]
  wire  _GEN_39226 = 6'h34 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39162; // @[rob.scala 181:{35,35}]
  wire  _GEN_39227 = 6'h35 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39163; // @[rob.scala 181:{35,35}]
  wire  _GEN_39228 = 6'h36 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39164; // @[rob.scala 181:{35,35}]
  wire  _GEN_39229 = 6'h37 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39165; // @[rob.scala 181:{35,35}]
  wire  _GEN_39230 = 6'h38 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39166; // @[rob.scala 181:{35,35}]
  wire  _GEN_39231 = 6'h39 == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39167; // @[rob.scala 181:{35,35}]
  wire  _GEN_39232 = 6'h3a == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39168; // @[rob.scala 181:{35,35}]
  wire  _GEN_39233 = 6'h3b == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39169; // @[rob.scala 181:{35,35}]
  wire  _GEN_39234 = 6'h3c == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39170; // @[rob.scala 181:{35,35}]
  wire  _GEN_39235 = 6'h3d == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39171; // @[rob.scala 181:{35,35}]
  wire  _GEN_39236 = 6'h3e == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39172; // @[rob.scala 181:{35,35}]
  wire  _GEN_39237 = 6'h3f == _next_can_commit_1_T_1[5:0] ? 1'h0 : _GEN_39173; // @[rob.scala 181:{35,35}]
  wire  _GEN_39302 = next_will_commit_0 ? _GEN_39110 : _GEN_36934; // @[rob.scala 183:38]
  wire  _GEN_39303 = next_will_commit_0 ? _GEN_39111 : _GEN_36935; // @[rob.scala 183:38]
  wire  _GEN_39304 = next_will_commit_0 ? _GEN_39112 : _GEN_36936; // @[rob.scala 183:38]
  wire  _GEN_39305 = next_will_commit_0 ? _GEN_39113 : _GEN_36937; // @[rob.scala 183:38]
  wire  _GEN_39306 = next_will_commit_0 ? _GEN_39114 : _GEN_36938; // @[rob.scala 183:38]
  wire  _GEN_39307 = next_will_commit_0 ? _GEN_39115 : _GEN_36939; // @[rob.scala 183:38]
  wire  _GEN_39308 = next_will_commit_0 ? _GEN_39116 : _GEN_36940; // @[rob.scala 183:38]
  wire  _GEN_39309 = next_will_commit_0 ? _GEN_39117 : _GEN_36941; // @[rob.scala 183:38]
  wire  _GEN_39310 = next_will_commit_0 ? _GEN_39118 : _GEN_36942; // @[rob.scala 183:38]
  wire  _GEN_39311 = next_will_commit_0 ? _GEN_39119 : _GEN_36943; // @[rob.scala 183:38]
  wire  _GEN_39312 = next_will_commit_0 ? _GEN_39120 : _GEN_36944; // @[rob.scala 183:38]
  wire  _GEN_39313 = next_will_commit_0 ? _GEN_39121 : _GEN_36945; // @[rob.scala 183:38]
  wire  _GEN_39314 = next_will_commit_0 ? _GEN_39122 : _GEN_36946; // @[rob.scala 183:38]
  wire  _GEN_39315 = next_will_commit_0 ? _GEN_39123 : _GEN_36947; // @[rob.scala 183:38]
  wire  _GEN_39316 = next_will_commit_0 ? _GEN_39124 : _GEN_36948; // @[rob.scala 183:38]
  wire  _GEN_39317 = next_will_commit_0 ? _GEN_39125 : _GEN_36949; // @[rob.scala 183:38]
  wire  _GEN_39318 = next_will_commit_0 ? _GEN_39126 : _GEN_36950; // @[rob.scala 183:38]
  wire  _GEN_39319 = next_will_commit_0 ? _GEN_39127 : _GEN_36951; // @[rob.scala 183:38]
  wire  _GEN_39320 = next_will_commit_0 ? _GEN_39128 : _GEN_36952; // @[rob.scala 183:38]
  wire  _GEN_39321 = next_will_commit_0 ? _GEN_39129 : _GEN_36953; // @[rob.scala 183:38]
  wire  _GEN_39322 = next_will_commit_0 ? _GEN_39130 : _GEN_36954; // @[rob.scala 183:38]
  wire  _GEN_39323 = next_will_commit_0 ? _GEN_39131 : _GEN_36955; // @[rob.scala 183:38]
  wire  _GEN_39324 = next_will_commit_0 ? _GEN_39132 : _GEN_36956; // @[rob.scala 183:38]
  wire  _GEN_39325 = next_will_commit_0 ? _GEN_39133 : _GEN_36957; // @[rob.scala 183:38]
  wire  _GEN_39326 = next_will_commit_0 ? _GEN_39134 : _GEN_36958; // @[rob.scala 183:38]
  wire  _GEN_39327 = next_will_commit_0 ? _GEN_39135 : _GEN_36959; // @[rob.scala 183:38]
  wire  _GEN_39328 = next_will_commit_0 ? _GEN_39136 : _GEN_36960; // @[rob.scala 183:38]
  wire  _GEN_39329 = next_will_commit_0 ? _GEN_39137 : _GEN_36961; // @[rob.scala 183:38]
  wire  _GEN_39330 = next_will_commit_0 ? _GEN_39138 : _GEN_36962; // @[rob.scala 183:38]
  wire  _GEN_39331 = next_will_commit_0 ? _GEN_39139 : _GEN_36963; // @[rob.scala 183:38]
  wire  _GEN_39332 = next_will_commit_0 ? _GEN_39140 : _GEN_36964; // @[rob.scala 183:38]
  wire  _GEN_39333 = next_will_commit_0 ? _GEN_39141 : _GEN_36965; // @[rob.scala 183:38]
  wire  _GEN_39334 = next_will_commit_0 ? _GEN_39142 : _GEN_36966; // @[rob.scala 183:38]
  wire  _GEN_39335 = next_will_commit_0 ? _GEN_39143 : _GEN_36967; // @[rob.scala 183:38]
  wire  _GEN_39336 = next_will_commit_0 ? _GEN_39144 : _GEN_36968; // @[rob.scala 183:38]
  wire  _GEN_39337 = next_will_commit_0 ? _GEN_39145 : _GEN_36969; // @[rob.scala 183:38]
  wire  _GEN_39338 = next_will_commit_0 ? _GEN_39146 : _GEN_36970; // @[rob.scala 183:38]
  wire  _GEN_39339 = next_will_commit_0 ? _GEN_39147 : _GEN_36971; // @[rob.scala 183:38]
  wire  _GEN_39340 = next_will_commit_0 ? _GEN_39148 : _GEN_36972; // @[rob.scala 183:38]
  wire  _GEN_39341 = next_will_commit_0 ? _GEN_39149 : _GEN_36973; // @[rob.scala 183:38]
  wire  _GEN_39342 = next_will_commit_0 ? _GEN_39150 : _GEN_36974; // @[rob.scala 183:38]
  wire  _GEN_39343 = next_will_commit_0 ? _GEN_39151 : _GEN_36975; // @[rob.scala 183:38]
  wire  _GEN_39344 = next_will_commit_0 ? _GEN_39152 : _GEN_36976; // @[rob.scala 183:38]
  wire  _GEN_39345 = next_will_commit_0 ? _GEN_39153 : _GEN_36977; // @[rob.scala 183:38]
  wire  _GEN_39346 = next_will_commit_0 ? _GEN_39154 : _GEN_36978; // @[rob.scala 183:38]
  wire  _GEN_39347 = next_will_commit_0 ? _GEN_39155 : _GEN_36979; // @[rob.scala 183:38]
  wire  _GEN_39348 = next_will_commit_0 ? _GEN_39156 : _GEN_36980; // @[rob.scala 183:38]
  wire  _GEN_39349 = next_will_commit_0 ? _GEN_39157 : _GEN_36981; // @[rob.scala 183:38]
  wire  _GEN_39350 = next_will_commit_0 ? _GEN_39158 : _GEN_36982; // @[rob.scala 183:38]
  wire  _GEN_39351 = next_will_commit_0 ? _GEN_39159 : _GEN_36983; // @[rob.scala 183:38]
  wire  _GEN_39352 = next_will_commit_0 ? _GEN_39160 : _GEN_36984; // @[rob.scala 183:38]
  wire  _GEN_39353 = next_will_commit_0 ? _GEN_39161 : _GEN_36985; // @[rob.scala 183:38]
  wire  _GEN_39354 = next_will_commit_0 ? _GEN_39162 : _GEN_36986; // @[rob.scala 183:38]
  wire  _GEN_39355 = next_will_commit_0 ? _GEN_39163 : _GEN_36987; // @[rob.scala 183:38]
  wire  _GEN_39356 = next_will_commit_0 ? _GEN_39164 : _GEN_36988; // @[rob.scala 183:38]
  wire  _GEN_39357 = next_will_commit_0 ? _GEN_39165 : _GEN_36989; // @[rob.scala 183:38]
  wire  _GEN_39358 = next_will_commit_0 ? _GEN_39166 : _GEN_36990; // @[rob.scala 183:38]
  wire  _GEN_39359 = next_will_commit_0 ? _GEN_39167 : _GEN_36991; // @[rob.scala 183:38]
  wire  _GEN_39360 = next_will_commit_0 ? _GEN_39168 : _GEN_36992; // @[rob.scala 183:38]
  wire  _GEN_39361 = next_will_commit_0 ? _GEN_39169 : _GEN_36993; // @[rob.scala 183:38]
  wire  _GEN_39362 = next_will_commit_0 ? _GEN_39170 : _GEN_36994; // @[rob.scala 183:38]
  wire  _GEN_39363 = next_will_commit_0 ? _GEN_39171 : _GEN_36995; // @[rob.scala 183:38]
  wire  _GEN_39364 = next_will_commit_0 ? _GEN_39172 : _GEN_36996; // @[rob.scala 183:38]
  wire  _GEN_39365 = next_will_commit_0 ? _GEN_39173 : _GEN_36997; // @[rob.scala 183:38]
  wire [6:0] _GEN_39366 = next_will_commit_0 ? _next_can_commit_1_T_1 : _GEN_30405; // @[rob.scala 183:38 185:20]
  wire  _GEN_39367 = _T_26 ? _GEN_39174 : _GEN_39302; // @[rob.scala 179:55]
  wire  _GEN_39368 = _T_26 ? _GEN_39175 : _GEN_39303; // @[rob.scala 179:55]
  wire  _GEN_39369 = _T_26 ? _GEN_39176 : _GEN_39304; // @[rob.scala 179:55]
  wire  _GEN_39370 = _T_26 ? _GEN_39177 : _GEN_39305; // @[rob.scala 179:55]
  wire  _GEN_39371 = _T_26 ? _GEN_39178 : _GEN_39306; // @[rob.scala 179:55]
  wire  _GEN_39372 = _T_26 ? _GEN_39179 : _GEN_39307; // @[rob.scala 179:55]
  wire  _GEN_39373 = _T_26 ? _GEN_39180 : _GEN_39308; // @[rob.scala 179:55]
  wire  _GEN_39374 = _T_26 ? _GEN_39181 : _GEN_39309; // @[rob.scala 179:55]
  wire  _GEN_39375 = _T_26 ? _GEN_39182 : _GEN_39310; // @[rob.scala 179:55]
  wire  _GEN_39376 = _T_26 ? _GEN_39183 : _GEN_39311; // @[rob.scala 179:55]
  wire  _GEN_39377 = _T_26 ? _GEN_39184 : _GEN_39312; // @[rob.scala 179:55]
  wire  _GEN_39378 = _T_26 ? _GEN_39185 : _GEN_39313; // @[rob.scala 179:55]
  wire  _GEN_39379 = _T_26 ? _GEN_39186 : _GEN_39314; // @[rob.scala 179:55]
  wire  _GEN_39380 = _T_26 ? _GEN_39187 : _GEN_39315; // @[rob.scala 179:55]
  wire  _GEN_39381 = _T_26 ? _GEN_39188 : _GEN_39316; // @[rob.scala 179:55]
  wire  _GEN_39382 = _T_26 ? _GEN_39189 : _GEN_39317; // @[rob.scala 179:55]
  wire  _GEN_39383 = _T_26 ? _GEN_39190 : _GEN_39318; // @[rob.scala 179:55]
  wire  _GEN_39384 = _T_26 ? _GEN_39191 : _GEN_39319; // @[rob.scala 179:55]
  wire  _GEN_39385 = _T_26 ? _GEN_39192 : _GEN_39320; // @[rob.scala 179:55]
  wire  _GEN_39386 = _T_26 ? _GEN_39193 : _GEN_39321; // @[rob.scala 179:55]
  wire  _GEN_39387 = _T_26 ? _GEN_39194 : _GEN_39322; // @[rob.scala 179:55]
  wire  _GEN_39388 = _T_26 ? _GEN_39195 : _GEN_39323; // @[rob.scala 179:55]
  wire  _GEN_39389 = _T_26 ? _GEN_39196 : _GEN_39324; // @[rob.scala 179:55]
  wire  _GEN_39390 = _T_26 ? _GEN_39197 : _GEN_39325; // @[rob.scala 179:55]
  wire  _GEN_39391 = _T_26 ? _GEN_39198 : _GEN_39326; // @[rob.scala 179:55]
  wire  _GEN_39392 = _T_26 ? _GEN_39199 : _GEN_39327; // @[rob.scala 179:55]
  wire  _GEN_39393 = _T_26 ? _GEN_39200 : _GEN_39328; // @[rob.scala 179:55]
  wire  _GEN_39394 = _T_26 ? _GEN_39201 : _GEN_39329; // @[rob.scala 179:55]
  wire  _GEN_39395 = _T_26 ? _GEN_39202 : _GEN_39330; // @[rob.scala 179:55]
  wire  _GEN_39396 = _T_26 ? _GEN_39203 : _GEN_39331; // @[rob.scala 179:55]
  wire  _GEN_39397 = _T_26 ? _GEN_39204 : _GEN_39332; // @[rob.scala 179:55]
  wire  _GEN_39398 = _T_26 ? _GEN_39205 : _GEN_39333; // @[rob.scala 179:55]
  wire  _GEN_39399 = _T_26 ? _GEN_39206 : _GEN_39334; // @[rob.scala 179:55]
  wire  _GEN_39400 = _T_26 ? _GEN_39207 : _GEN_39335; // @[rob.scala 179:55]
  wire  _GEN_39401 = _T_26 ? _GEN_39208 : _GEN_39336; // @[rob.scala 179:55]
  wire  _GEN_39402 = _T_26 ? _GEN_39209 : _GEN_39337; // @[rob.scala 179:55]
  wire  _GEN_39403 = _T_26 ? _GEN_39210 : _GEN_39338; // @[rob.scala 179:55]
  wire  _GEN_39404 = _T_26 ? _GEN_39211 : _GEN_39339; // @[rob.scala 179:55]
  wire  _GEN_39405 = _T_26 ? _GEN_39212 : _GEN_39340; // @[rob.scala 179:55]
  wire  _GEN_39406 = _T_26 ? _GEN_39213 : _GEN_39341; // @[rob.scala 179:55]
  wire  _GEN_39407 = _T_26 ? _GEN_39214 : _GEN_39342; // @[rob.scala 179:55]
  wire  _GEN_39408 = _T_26 ? _GEN_39215 : _GEN_39343; // @[rob.scala 179:55]
  wire  _GEN_39409 = _T_26 ? _GEN_39216 : _GEN_39344; // @[rob.scala 179:55]
  wire  _GEN_39410 = _T_26 ? _GEN_39217 : _GEN_39345; // @[rob.scala 179:55]
  wire  _GEN_39411 = _T_26 ? _GEN_39218 : _GEN_39346; // @[rob.scala 179:55]
  wire  _GEN_39412 = _T_26 ? _GEN_39219 : _GEN_39347; // @[rob.scala 179:55]
  wire  _GEN_39413 = _T_26 ? _GEN_39220 : _GEN_39348; // @[rob.scala 179:55]
  wire  _GEN_39414 = _T_26 ? _GEN_39221 : _GEN_39349; // @[rob.scala 179:55]
  wire  _GEN_39415 = _T_26 ? _GEN_39222 : _GEN_39350; // @[rob.scala 179:55]
  wire  _GEN_39416 = _T_26 ? _GEN_39223 : _GEN_39351; // @[rob.scala 179:55]
  wire  _GEN_39417 = _T_26 ? _GEN_39224 : _GEN_39352; // @[rob.scala 179:55]
  wire  _GEN_39418 = _T_26 ? _GEN_39225 : _GEN_39353; // @[rob.scala 179:55]
  wire  _GEN_39419 = _T_26 ? _GEN_39226 : _GEN_39354; // @[rob.scala 179:55]
  wire  _GEN_39420 = _T_26 ? _GEN_39227 : _GEN_39355; // @[rob.scala 179:55]
  wire  _GEN_39421 = _T_26 ? _GEN_39228 : _GEN_39356; // @[rob.scala 179:55]
  wire  _GEN_39422 = _T_26 ? _GEN_39229 : _GEN_39357; // @[rob.scala 179:55]
  wire  _GEN_39423 = _T_26 ? _GEN_39230 : _GEN_39358; // @[rob.scala 179:55]
  wire  _GEN_39424 = _T_26 ? _GEN_39231 : _GEN_39359; // @[rob.scala 179:55]
  wire  _GEN_39425 = _T_26 ? _GEN_39232 : _GEN_39360; // @[rob.scala 179:55]
  wire  _GEN_39426 = _T_26 ? _GEN_39233 : _GEN_39361; // @[rob.scala 179:55]
  wire  _GEN_39427 = _T_26 ? _GEN_39234 : _GEN_39362; // @[rob.scala 179:55]
  wire  _GEN_39428 = _T_26 ? _GEN_39235 : _GEN_39363; // @[rob.scala 179:55]
  wire  _GEN_39429 = _T_26 ? _GEN_39236 : _GEN_39364; // @[rob.scala 179:55]
  wire  _GEN_39430 = _T_26 ? _GEN_39237 : _GEN_39365; // @[rob.scala 179:55]
  wire  _GEN_39432 = _next_will_commit_0_T_6 ? _GEN_39367 : _GEN_30212; // @[rob.scala 164:36]
  wire  _GEN_39433 = _next_will_commit_0_T_6 ? _GEN_39368 : _GEN_30213; // @[rob.scala 164:36]
  wire  _GEN_39434 = _next_will_commit_0_T_6 ? _GEN_39369 : _GEN_30214; // @[rob.scala 164:36]
  wire  _GEN_39435 = _next_will_commit_0_T_6 ? _GEN_39370 : _GEN_30215; // @[rob.scala 164:36]
  wire  _GEN_39436 = _next_will_commit_0_T_6 ? _GEN_39371 : _GEN_30216; // @[rob.scala 164:36]
  wire  _GEN_39437 = _next_will_commit_0_T_6 ? _GEN_39372 : _GEN_30217; // @[rob.scala 164:36]
  wire  _GEN_39438 = _next_will_commit_0_T_6 ? _GEN_39373 : _GEN_30218; // @[rob.scala 164:36]
  wire  _GEN_39439 = _next_will_commit_0_T_6 ? _GEN_39374 : _GEN_30219; // @[rob.scala 164:36]
  wire  _GEN_39440 = _next_will_commit_0_T_6 ? _GEN_39375 : _GEN_30220; // @[rob.scala 164:36]
  wire  _GEN_39441 = _next_will_commit_0_T_6 ? _GEN_39376 : _GEN_30221; // @[rob.scala 164:36]
  wire  _GEN_39442 = _next_will_commit_0_T_6 ? _GEN_39377 : _GEN_30222; // @[rob.scala 164:36]
  wire  _GEN_39443 = _next_will_commit_0_T_6 ? _GEN_39378 : _GEN_30223; // @[rob.scala 164:36]
  wire  _GEN_39444 = _next_will_commit_0_T_6 ? _GEN_39379 : _GEN_30224; // @[rob.scala 164:36]
  wire  _GEN_39445 = _next_will_commit_0_T_6 ? _GEN_39380 : _GEN_30225; // @[rob.scala 164:36]
  wire  _GEN_39446 = _next_will_commit_0_T_6 ? _GEN_39381 : _GEN_30226; // @[rob.scala 164:36]
  wire  _GEN_39447 = _next_will_commit_0_T_6 ? _GEN_39382 : _GEN_30227; // @[rob.scala 164:36]
  wire  _GEN_39448 = _next_will_commit_0_T_6 ? _GEN_39383 : _GEN_30228; // @[rob.scala 164:36]
  wire  _GEN_39449 = _next_will_commit_0_T_6 ? _GEN_39384 : _GEN_30229; // @[rob.scala 164:36]
  wire  _GEN_39450 = _next_will_commit_0_T_6 ? _GEN_39385 : _GEN_30230; // @[rob.scala 164:36]
  wire  _GEN_39451 = _next_will_commit_0_T_6 ? _GEN_39386 : _GEN_30231; // @[rob.scala 164:36]
  wire  _GEN_39452 = _next_will_commit_0_T_6 ? _GEN_39387 : _GEN_30232; // @[rob.scala 164:36]
  wire  _GEN_39453 = _next_will_commit_0_T_6 ? _GEN_39388 : _GEN_30233; // @[rob.scala 164:36]
  wire  _GEN_39454 = _next_will_commit_0_T_6 ? _GEN_39389 : _GEN_30234; // @[rob.scala 164:36]
  wire  _GEN_39455 = _next_will_commit_0_T_6 ? _GEN_39390 : _GEN_30235; // @[rob.scala 164:36]
  wire  _GEN_39456 = _next_will_commit_0_T_6 ? _GEN_39391 : _GEN_30236; // @[rob.scala 164:36]
  wire  _GEN_39457 = _next_will_commit_0_T_6 ? _GEN_39392 : _GEN_30237; // @[rob.scala 164:36]
  wire  _GEN_39458 = _next_will_commit_0_T_6 ? _GEN_39393 : _GEN_30238; // @[rob.scala 164:36]
  wire  _GEN_39459 = _next_will_commit_0_T_6 ? _GEN_39394 : _GEN_30239; // @[rob.scala 164:36]
  wire  _GEN_39460 = _next_will_commit_0_T_6 ? _GEN_39395 : _GEN_30240; // @[rob.scala 164:36]
  wire  _GEN_39461 = _next_will_commit_0_T_6 ? _GEN_39396 : _GEN_30241; // @[rob.scala 164:36]
  wire  _GEN_39462 = _next_will_commit_0_T_6 ? _GEN_39397 : _GEN_30242; // @[rob.scala 164:36]
  wire  _GEN_39463 = _next_will_commit_0_T_6 ? _GEN_39398 : _GEN_30243; // @[rob.scala 164:36]
  wire  _GEN_39464 = _next_will_commit_0_T_6 ? _GEN_39399 : _GEN_30244; // @[rob.scala 164:36]
  wire  _GEN_39465 = _next_will_commit_0_T_6 ? _GEN_39400 : _GEN_30245; // @[rob.scala 164:36]
  wire  _GEN_39466 = _next_will_commit_0_T_6 ? _GEN_39401 : _GEN_30246; // @[rob.scala 164:36]
  wire  _GEN_39467 = _next_will_commit_0_T_6 ? _GEN_39402 : _GEN_30247; // @[rob.scala 164:36]
  wire  _GEN_39468 = _next_will_commit_0_T_6 ? _GEN_39403 : _GEN_30248; // @[rob.scala 164:36]
  wire  _GEN_39469 = _next_will_commit_0_T_6 ? _GEN_39404 : _GEN_30249; // @[rob.scala 164:36]
  wire  _GEN_39470 = _next_will_commit_0_T_6 ? _GEN_39405 : _GEN_30250; // @[rob.scala 164:36]
  wire  _GEN_39471 = _next_will_commit_0_T_6 ? _GEN_39406 : _GEN_30251; // @[rob.scala 164:36]
  wire  _GEN_39472 = _next_will_commit_0_T_6 ? _GEN_39407 : _GEN_30252; // @[rob.scala 164:36]
  wire  _GEN_39473 = _next_will_commit_0_T_6 ? _GEN_39408 : _GEN_30253; // @[rob.scala 164:36]
  wire  _GEN_39474 = _next_will_commit_0_T_6 ? _GEN_39409 : _GEN_30254; // @[rob.scala 164:36]
  wire  _GEN_39475 = _next_will_commit_0_T_6 ? _GEN_39410 : _GEN_30255; // @[rob.scala 164:36]
  wire  _GEN_39476 = _next_will_commit_0_T_6 ? _GEN_39411 : _GEN_30256; // @[rob.scala 164:36]
  wire  _GEN_39477 = _next_will_commit_0_T_6 ? _GEN_39412 : _GEN_30257; // @[rob.scala 164:36]
  wire  _GEN_39478 = _next_will_commit_0_T_6 ? _GEN_39413 : _GEN_30258; // @[rob.scala 164:36]
  wire  _GEN_39479 = _next_will_commit_0_T_6 ? _GEN_39414 : _GEN_30259; // @[rob.scala 164:36]
  wire  _GEN_39480 = _next_will_commit_0_T_6 ? _GEN_39415 : _GEN_30260; // @[rob.scala 164:36]
  wire  _GEN_39481 = _next_will_commit_0_T_6 ? _GEN_39416 : _GEN_30261; // @[rob.scala 164:36]
  wire  _GEN_39482 = _next_will_commit_0_T_6 ? _GEN_39417 : _GEN_30262; // @[rob.scala 164:36]
  wire  _GEN_39483 = _next_will_commit_0_T_6 ? _GEN_39418 : _GEN_30263; // @[rob.scala 164:36]
  wire  _GEN_39484 = _next_will_commit_0_T_6 ? _GEN_39419 : _GEN_30264; // @[rob.scala 164:36]
  wire  _GEN_39485 = _next_will_commit_0_T_6 ? _GEN_39420 : _GEN_30265; // @[rob.scala 164:36]
  wire  _GEN_39486 = _next_will_commit_0_T_6 ? _GEN_39421 : _GEN_30266; // @[rob.scala 164:36]
  wire  _GEN_39487 = _next_will_commit_0_T_6 ? _GEN_39422 : _GEN_30267; // @[rob.scala 164:36]
  wire  _GEN_39488 = _next_will_commit_0_T_6 ? _GEN_39423 : _GEN_30268; // @[rob.scala 164:36]
  wire  _GEN_39489 = _next_will_commit_0_T_6 ? _GEN_39424 : _GEN_30269; // @[rob.scala 164:36]
  wire  _GEN_39490 = _next_will_commit_0_T_6 ? _GEN_39425 : _GEN_30270; // @[rob.scala 164:36]
  wire  _GEN_39491 = _next_will_commit_0_T_6 ? _GEN_39426 : _GEN_30271; // @[rob.scala 164:36]
  wire  _GEN_39492 = _next_will_commit_0_T_6 ? _GEN_39427 : _GEN_30272; // @[rob.scala 164:36]
  wire  _GEN_39493 = _next_will_commit_0_T_6 ? _GEN_39428 : _GEN_30273; // @[rob.scala 164:36]
  wire  _GEN_39494 = _next_will_commit_0_T_6 ? _GEN_39429 : _GEN_30274; // @[rob.scala 164:36]
  wire  _GEN_39495 = _next_will_commit_0_T_6 ? _GEN_39430 : _GEN_30275; // @[rob.scala 164:36]
  wire [6:0] _allocate_ptr_T_5 = allocate_ptr - this_num_to_roll_back; // @[rob.scala 190:36]
  assign io_o_full = _is_full_T_1 == commit_ptr | _is_full_T_4 == commit_ptr; // @[rob.scala 208:52]
  assign io_o_rob_allocation_ress_0_rob_idx = allocate_ptr; // @[rob.scala 120:43]
  assign io_o_rob_allocation_ress_1_rob_idx = allocate_ptr + 7'h1; // @[rob.scala 121:58]
  assign io_o_rollback_packs_0_valid = next_rob_state == 2'h2; // @[rob.scala 114:53]
  assign io_o_rollback_packs_0_uop_phy_dst = 6'h3f == _next_rob_state_T_10[5:0] ? rob_uop_63_phy_dst : _GEN_5310; // @[rob.scala 117:{33,33}]
  assign io_o_rollback_packs_0_uop_stale_dst = 6'h3f == _next_rob_state_T_10[5:0] ? rob_uop_63_stale_dst : _GEN_5374; // @[rob.scala 117:{33,33}]
  assign io_o_rollback_packs_0_uop_arch_dst = 6'h3f == _next_rob_state_T_10[5:0] ? rob_uop_63_arch_dst : _GEN_5438; // @[rob.scala 117:{33,33}]
  assign io_o_rollback_packs_1_valid = this_num_to_roll_back == 7'h2 & _this_num_to_roll_back_T; // @[rob.scala 115:71]
  assign io_o_rollback_packs_1_uop_phy_dst = 6'h3f == _next_rob_state_T_13[5:0] ? rob_uop_63_phy_dst : _GEN_7294; // @[rob.scala 118:{33,33}]
  assign io_o_rollback_packs_1_uop_stale_dst = 6'h3f == _next_rob_state_T_13[5:0] ? rob_uop_63_stale_dst : _GEN_7358; // @[rob.scala 118:{33,33}]
  assign io_o_rollback_packs_1_uop_arch_dst = 6'h3f == _next_rob_state_T_13[5:0] ? rob_uop_63_arch_dst : _GEN_7422; // @[rob.scala 118:{33,33}]
  assign io_o_commit_packs_0_valid = next_will_commit_0 & _next_will_commit_0_T_7; // @[rob.scala 106:59]
  assign io_o_commit_packs_0_uop_pc = 6'h3f == commit_ptr[5:0] ? rob_uop_63_pc : _GEN_830; // @[rob.scala 108:{32,32}]
  assign io_o_commit_packs_0_uop_inst = 6'h3f == commit_ptr[5:0] ? rob_uop_63_inst : _GEN_894; // @[rob.scala 108:{32,32}]
  assign io_o_commit_packs_0_uop_func_code = 6'h3f == commit_ptr[5:0] ? rob_uop_63_func_code : _GEN_382; // @[rob.scala 108:{32,32}]
  assign io_o_commit_packs_0_uop_phy_dst = 6'h3f == commit_ptr[5:0] ? rob_uop_63_phy_dst : _GEN_1342; // @[rob.scala 108:{32,32}]
  assign io_o_commit_packs_0_uop_stale_dst = 6'h3f == commit_ptr[5:0] ? rob_uop_63_stale_dst : _GEN_1406; // @[rob.scala 108:{32,32}]
  assign io_o_commit_packs_0_uop_arch_dst = 6'h3f == commit_ptr[5:0] ? rob_uop_63_arch_dst : _GEN_1470; // @[rob.scala 108:{32,32}]
  assign io_o_commit_packs_0_uop_dst_value = 6'h3f == commit_ptr[5:0] ? rob_uop_63_dst_value : _GEN_2174; // @[rob.scala 108:{32,32}]
  assign io_o_commit_packs_0_uop_src1_value = 6'h3f == commit_ptr[5:0] ? rob_uop_63_src1_value : _GEN_2238; // @[rob.scala 108:{32,32}]
  assign io_o_commit_packs_0_uop_alu_sel = 6'h3f == commit_ptr[5:0] ? rob_uop_63_alu_sel : _GEN_446; // @[rob.scala 108:{32,32}]
  assign io_o_commit_packs_1_valid = next_will_commit_1 & next_will_commit_0 & _next_will_commit_0_T_7; // @[rob.scala 107:82]
  assign io_o_commit_packs_1_uop_inst = 6'h3f == _next_can_commit_1_T_1[5:0] ? rob_uop_63_inst : _GEN_2878; // @[rob.scala 109:{32,32}]
  assign io_o_commit_packs_1_uop_func_code = 6'h3f == _next_can_commit_1_T_1[5:0] ? rob_uop_63_func_code : _GEN_2942; // @[rob.scala 109:{32,32}]
  assign io_o_commit_packs_1_uop_phy_dst = 6'h3f == _next_can_commit_1_T_1[5:0] ? rob_uop_63_phy_dst : _GEN_3326; // @[rob.scala 109:{32,32}]
  assign io_o_commit_packs_1_uop_stale_dst = 6'h3f == _next_can_commit_1_T_1[5:0] ? rob_uop_63_stale_dst : _GEN_3390; // @[rob.scala 109:{32,32}]
  assign io_o_commit_packs_1_uop_arch_dst = 6'h3f == _next_can_commit_1_T_1[5:0] ? rob_uop_63_arch_dst : _GEN_3454; // @[rob.scala 109:{32,32}]
  assign io_o_commit_packs_1_uop_dst_value = 6'h3f == _next_can_commit_1_T_1[5:0] ? rob_uop_63_dst_value : _GEN_4158; // @[rob.scala 109:{32,32}]
  assign io_o_commit_packs_1_uop_src1_value = 6'h3f == _next_can_commit_1_T_1[5:0] ? rob_uop_63_src1_value : _GEN_4222; // @[rob.scala 109:{32,32}]
  assign io_o_commit_packs_1_uop_alu_sel = 6'h3f == _next_can_commit_1_T_1[5:0] ? rob_uop_63_alu_sel : _GEN_4542; // @[rob.scala 109:{32,32}]
  assign io_o_rob_head = commit_ptr; // @[rob.scala 78:19]
  assign io_o_exception = 1'h0; // @[rob.scala 205:{47,47}]
  always @(posedge clock) begin
    if (reset) begin // @[rob.scala 46:29]
      commit_ptr <= 7'h0; // @[rob.scala 46:29]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      commit_ptr <= 7'h0; // @[rob.scala 198:20]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (_T_26) begin // @[rob.scala 179:55]
        commit_ptr <= _commit_ptr_T_1; // @[rob.scala 182:20]
      end else begin
        commit_ptr <= _GEN_39366;
      end
    end else if (_next_will_commit_0_T_5) begin // @[rob.scala 123:38]
      commit_ptr <= _GEN_28227;
    end
    if (reset) begin // @[rob.scala 47:31]
      allocate_ptr <= 7'h0; // @[rob.scala 47:31]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      allocate_ptr <= 7'h0; // @[rob.scala 197:22]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      allocate_ptr <= _allocate_ptr_T_5; // @[rob.scala 190:20]
    end else if (_next_will_commit_0_T_5) begin // @[rob.scala 123:38]
      allocate_ptr <= _GEN_19201;
    end
    if (reset) begin // @[rob.scala 53:28]
      rob_state <= 2'h1; // @[rob.scala 53:28]
    end else if (io_o_exception | io_i_interrupt | last_pc_redirect) begin // @[rob.scala 214:24]
      rob_state <= 2'h0;
    end else if (_next_rob_state_T_2) begin // @[Mux.scala 101:16]
      rob_state <= 2'h1;
    end else if (_next_rob_state_T_4) begin // @[Mux.scala 101:16]
      rob_state <= 2'h3;
    end else begin
      rob_state <= _next_rob_state_T_21;
    end
    last_pc_redirect <= io_i_csr_pc_redirect; // @[rob.scala 56:22]
    if (reset) begin // @[rob.scala 89:30]
      will_commit_0 <= 1'h0; // @[rob.scala 89:30]
    end else begin
      will_commit_0 <= next_will_commit_0; // @[rob.scala 91:17]
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_0 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_0 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h0 == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_0 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_0 <= _GEN_39432;
      end
    end else begin
      rob_valid_0 <= _GEN_39432;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_1 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_1 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h1 == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_1 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_1 <= _GEN_39433;
      end
    end else begin
      rob_valid_1 <= _GEN_39433;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_2 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_2 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h2 == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_2 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_2 <= _GEN_39434;
      end
    end else begin
      rob_valid_2 <= _GEN_39434;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_3 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_3 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h3 == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_3 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_3 <= _GEN_39435;
      end
    end else begin
      rob_valid_3 <= _GEN_39435;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_4 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_4 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h4 == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_4 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_4 <= _GEN_39436;
      end
    end else begin
      rob_valid_4 <= _GEN_39436;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_5 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_5 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h5 == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_5 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_5 <= _GEN_39437;
      end
    end else begin
      rob_valid_5 <= _GEN_39437;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_6 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_6 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h6 == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_6 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_6 <= _GEN_39438;
      end
    end else begin
      rob_valid_6 <= _GEN_39438;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_7 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_7 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h7 == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_7 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_7 <= _GEN_39439;
      end
    end else begin
      rob_valid_7 <= _GEN_39439;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_8 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_8 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h8 == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_8 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_8 <= _GEN_39440;
      end
    end else begin
      rob_valid_8 <= _GEN_39440;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_9 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_9 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h9 == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_9 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_9 <= _GEN_39441;
      end
    end else begin
      rob_valid_9 <= _GEN_39441;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_10 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_10 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'ha == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_10 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_10 <= _GEN_39442;
      end
    end else begin
      rob_valid_10 <= _GEN_39442;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_11 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_11 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'hb == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_11 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_11 <= _GEN_39443;
      end
    end else begin
      rob_valid_11 <= _GEN_39443;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_12 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_12 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'hc == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_12 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_12 <= _GEN_39444;
      end
    end else begin
      rob_valid_12 <= _GEN_39444;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_13 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_13 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'hd == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_13 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_13 <= _GEN_39445;
      end
    end else begin
      rob_valid_13 <= _GEN_39445;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_14 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_14 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'he == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_14 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_14 <= _GEN_39446;
      end
    end else begin
      rob_valid_14 <= _GEN_39446;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_15 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_15 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'hf == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_15 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_15 <= _GEN_39447;
      end
    end else begin
      rob_valid_15 <= _GEN_39447;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_16 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_16 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h10 == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_16 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_16 <= _GEN_39448;
      end
    end else begin
      rob_valid_16 <= _GEN_39448;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_17 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_17 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h11 == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_17 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_17 <= _GEN_39449;
      end
    end else begin
      rob_valid_17 <= _GEN_39449;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_18 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_18 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h12 == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_18 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_18 <= _GEN_39450;
      end
    end else begin
      rob_valid_18 <= _GEN_39450;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_19 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_19 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h13 == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_19 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_19 <= _GEN_39451;
      end
    end else begin
      rob_valid_19 <= _GEN_39451;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_20 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_20 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h14 == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_20 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_20 <= _GEN_39452;
      end
    end else begin
      rob_valid_20 <= _GEN_39452;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_21 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_21 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h15 == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_21 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_21 <= _GEN_39453;
      end
    end else begin
      rob_valid_21 <= _GEN_39453;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_22 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_22 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h16 == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_22 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_22 <= _GEN_39454;
      end
    end else begin
      rob_valid_22 <= _GEN_39454;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_23 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_23 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h17 == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_23 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_23 <= _GEN_39455;
      end
    end else begin
      rob_valid_23 <= _GEN_39455;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_24 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_24 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h18 == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_24 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_24 <= _GEN_39456;
      end
    end else begin
      rob_valid_24 <= _GEN_39456;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_25 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_25 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h19 == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_25 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_25 <= _GEN_39457;
      end
    end else begin
      rob_valid_25 <= _GEN_39457;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_26 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_26 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h1a == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_26 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_26 <= _GEN_39458;
      end
    end else begin
      rob_valid_26 <= _GEN_39458;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_27 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_27 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h1b == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_27 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_27 <= _GEN_39459;
      end
    end else begin
      rob_valid_27 <= _GEN_39459;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_28 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_28 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h1c == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_28 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_28 <= _GEN_39460;
      end
    end else begin
      rob_valid_28 <= _GEN_39460;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_29 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_29 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h1d == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_29 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_29 <= _GEN_39461;
      end
    end else begin
      rob_valid_29 <= _GEN_39461;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_30 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_30 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h1e == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_30 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_30 <= _GEN_39462;
      end
    end else begin
      rob_valid_30 <= _GEN_39462;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_31 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_31 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h1f == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_31 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_31 <= _GEN_39463;
      end
    end else begin
      rob_valid_31 <= _GEN_39463;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_32 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_32 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h20 == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_32 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_32 <= _GEN_39464;
      end
    end else begin
      rob_valid_32 <= _GEN_39464;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_33 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_33 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h21 == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_33 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_33 <= _GEN_39465;
      end
    end else begin
      rob_valid_33 <= _GEN_39465;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_34 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_34 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h22 == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_34 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_34 <= _GEN_39466;
      end
    end else begin
      rob_valid_34 <= _GEN_39466;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_35 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_35 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h23 == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_35 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_35 <= _GEN_39467;
      end
    end else begin
      rob_valid_35 <= _GEN_39467;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_36 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_36 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h24 == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_36 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_36 <= _GEN_39468;
      end
    end else begin
      rob_valid_36 <= _GEN_39468;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_37 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_37 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h25 == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_37 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_37 <= _GEN_39469;
      end
    end else begin
      rob_valid_37 <= _GEN_39469;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_38 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_38 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h26 == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_38 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_38 <= _GEN_39470;
      end
    end else begin
      rob_valid_38 <= _GEN_39470;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_39 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_39 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h27 == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_39 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_39 <= _GEN_39471;
      end
    end else begin
      rob_valid_39 <= _GEN_39471;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_40 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_40 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h28 == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_40 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_40 <= _GEN_39472;
      end
    end else begin
      rob_valid_40 <= _GEN_39472;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_41 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_41 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h29 == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_41 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_41 <= _GEN_39473;
      end
    end else begin
      rob_valid_41 <= _GEN_39473;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_42 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_42 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h2a == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_42 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_42 <= _GEN_39474;
      end
    end else begin
      rob_valid_42 <= _GEN_39474;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_43 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_43 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h2b == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_43 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_43 <= _GEN_39475;
      end
    end else begin
      rob_valid_43 <= _GEN_39475;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_44 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_44 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h2c == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_44 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_44 <= _GEN_39476;
      end
    end else begin
      rob_valid_44 <= _GEN_39476;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_45 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_45 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h2d == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_45 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_45 <= _GEN_39477;
      end
    end else begin
      rob_valid_45 <= _GEN_39477;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_46 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_46 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h2e == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_46 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_46 <= _GEN_39478;
      end
    end else begin
      rob_valid_46 <= _GEN_39478;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_47 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_47 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h2f == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_47 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_47 <= _GEN_39479;
      end
    end else begin
      rob_valid_47 <= _GEN_39479;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_48 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_48 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h30 == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_48 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_48 <= _GEN_39480;
      end
    end else begin
      rob_valid_48 <= _GEN_39480;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_49 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_49 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h31 == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_49 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_49 <= _GEN_39481;
      end
    end else begin
      rob_valid_49 <= _GEN_39481;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_50 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_50 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h32 == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_50 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_50 <= _GEN_39482;
      end
    end else begin
      rob_valid_50 <= _GEN_39482;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_51 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_51 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h33 == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_51 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_51 <= _GEN_39483;
      end
    end else begin
      rob_valid_51 <= _GEN_39483;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_52 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_52 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h34 == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_52 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_52 <= _GEN_39484;
      end
    end else begin
      rob_valid_52 <= _GEN_39484;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_53 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_53 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h35 == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_53 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_53 <= _GEN_39485;
      end
    end else begin
      rob_valid_53 <= _GEN_39485;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_54 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_54 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h36 == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_54 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_54 <= _GEN_39486;
      end
    end else begin
      rob_valid_54 <= _GEN_39486;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_55 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_55 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h37 == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_55 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_55 <= _GEN_39487;
      end
    end else begin
      rob_valid_55 <= _GEN_39487;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_56 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_56 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h38 == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_56 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_56 <= _GEN_39488;
      end
    end else begin
      rob_valid_56 <= _GEN_39488;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_57 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_57 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h39 == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_57 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_57 <= _GEN_39489;
      end
    end else begin
      rob_valid_57 <= _GEN_39489;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_58 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_58 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h3a == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_58 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_58 <= _GEN_39490;
      end
    end else begin
      rob_valid_58 <= _GEN_39490;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_59 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_59 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h3b == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_59 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_59 <= _GEN_39491;
      end
    end else begin
      rob_valid_59 <= _GEN_39491;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_60 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_60 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h3c == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_60 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_60 <= _GEN_39492;
      end
    end else begin
      rob_valid_60 <= _GEN_39492;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_61 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_61 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h3d == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_61 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_61 <= _GEN_39493;
      end
    end else begin
      rob_valid_61 <= _GEN_39493;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_62 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_62 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h3e == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_62 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_62 <= _GEN_39494;
      end
    end else begin
      rob_valid_62 <= _GEN_39494;
    end
    if (reset) begin // @[rob.scala 81:28]
      rob_valid_63 <= 1'h0; // @[rob.scala 81:28]
    end else if (next_rob_state == 2'h0) begin // @[rob.scala 193:37]
      rob_valid_63 <= 1'h0; // @[rob.scala 195:24]
    end else if (_this_num_to_roll_back_T) begin // @[rob.scala 188:40]
      if (6'h3f == allocate_ptr[5:0]) begin // @[rob.scala 191:31]
        rob_valid_63 <= 1'h0; // @[rob.scala 191:31]
      end else begin
        rob_valid_63 <= _GEN_39495;
      end
    end else begin
      rob_valid_63 <= _GEN_39495;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_0_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h0 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_0_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_0_pc <= _GEN_32710;
        end
      end else begin
        rob_uop_0_pc <= _GEN_32710;
      end
    end else begin
      rob_uop_0_pc <= _GEN_28292;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_0_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h0 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_0_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_0_inst <= _GEN_32774;
        end
      end else begin
        rob_uop_0_inst <= _GEN_32774;
      end
    end else begin
      rob_uop_0_inst <= _GEN_28356;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_0_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h0 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_0_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_0_func_code <= _GEN_32838;
        end
      end else begin
        rob_uop_0_func_code <= _GEN_32838;
      end
    end else begin
      rob_uop_0_func_code <= _GEN_28420;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_0_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h0 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_0_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_0_phy_dst <= _GEN_33222;
        end
      end else begin
        rob_uop_0_phy_dst <= _GEN_33222;
      end
    end else begin
      rob_uop_0_phy_dst <= _GEN_28804;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_0_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h0 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_0_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_0_stale_dst <= _GEN_33286;
        end
      end else begin
        rob_uop_0_stale_dst <= _GEN_33286;
      end
    end else begin
      rob_uop_0_stale_dst <= _GEN_28868;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_0_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h0 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_0_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_0_arch_dst <= _GEN_33350;
        end
      end else begin
        rob_uop_0_arch_dst <= _GEN_33350;
      end
    end else begin
      rob_uop_0_arch_dst <= _GEN_28932;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_0_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h0 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_0_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_0_dst_value <= _GEN_34054;
        end
      end else begin
        rob_uop_0_dst_value <= _GEN_34054;
      end
    end else begin
      rob_uop_0_dst_value <= _GEN_29636;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_0_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h0 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_0_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_0_src1_value <= _GEN_34118;
        end
      end else begin
        rob_uop_0_src1_value <= _GEN_34118;
      end
    end else begin
      rob_uop_0_src1_value <= _GEN_29700;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_0_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h0 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_0_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_0_alu_sel <= _GEN_34438;
        end
      end else begin
        rob_uop_0_alu_sel <= _GEN_34438;
      end
    end else begin
      rob_uop_0_alu_sel <= _GEN_30020;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_1_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_1_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_1_pc <= _GEN_32711;
        end
      end else begin
        rob_uop_1_pc <= _GEN_32711;
      end
    end else begin
      rob_uop_1_pc <= _GEN_28293;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_1_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_1_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_1_inst <= _GEN_32775;
        end
      end else begin
        rob_uop_1_inst <= _GEN_32775;
      end
    end else begin
      rob_uop_1_inst <= _GEN_28357;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_1_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_1_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_1_func_code <= _GEN_32839;
        end
      end else begin
        rob_uop_1_func_code <= _GEN_32839;
      end
    end else begin
      rob_uop_1_func_code <= _GEN_28421;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_1_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_1_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_1_phy_dst <= _GEN_33223;
        end
      end else begin
        rob_uop_1_phy_dst <= _GEN_33223;
      end
    end else begin
      rob_uop_1_phy_dst <= _GEN_28805;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_1_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_1_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_1_stale_dst <= _GEN_33287;
        end
      end else begin
        rob_uop_1_stale_dst <= _GEN_33287;
      end
    end else begin
      rob_uop_1_stale_dst <= _GEN_28869;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_1_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_1_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_1_arch_dst <= _GEN_33351;
        end
      end else begin
        rob_uop_1_arch_dst <= _GEN_33351;
      end
    end else begin
      rob_uop_1_arch_dst <= _GEN_28933;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_1_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_1_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_1_dst_value <= _GEN_34055;
        end
      end else begin
        rob_uop_1_dst_value <= _GEN_34055;
      end
    end else begin
      rob_uop_1_dst_value <= _GEN_29637;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_1_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_1_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_1_src1_value <= _GEN_34119;
        end
      end else begin
        rob_uop_1_src1_value <= _GEN_34119;
      end
    end else begin
      rob_uop_1_src1_value <= _GEN_29701;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_1_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_1_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_1_alu_sel <= _GEN_34439;
        end
      end else begin
        rob_uop_1_alu_sel <= _GEN_34439;
      end
    end else begin
      rob_uop_1_alu_sel <= _GEN_30021;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_2_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_2_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_2_pc <= _GEN_32712;
        end
      end else begin
        rob_uop_2_pc <= _GEN_32712;
      end
    end else begin
      rob_uop_2_pc <= _GEN_28294;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_2_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_2_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_2_inst <= _GEN_32776;
        end
      end else begin
        rob_uop_2_inst <= _GEN_32776;
      end
    end else begin
      rob_uop_2_inst <= _GEN_28358;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_2_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_2_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_2_func_code <= _GEN_32840;
        end
      end else begin
        rob_uop_2_func_code <= _GEN_32840;
      end
    end else begin
      rob_uop_2_func_code <= _GEN_28422;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_2_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_2_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_2_phy_dst <= _GEN_33224;
        end
      end else begin
        rob_uop_2_phy_dst <= _GEN_33224;
      end
    end else begin
      rob_uop_2_phy_dst <= _GEN_28806;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_2_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_2_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_2_stale_dst <= _GEN_33288;
        end
      end else begin
        rob_uop_2_stale_dst <= _GEN_33288;
      end
    end else begin
      rob_uop_2_stale_dst <= _GEN_28870;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_2_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_2_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_2_arch_dst <= _GEN_33352;
        end
      end else begin
        rob_uop_2_arch_dst <= _GEN_33352;
      end
    end else begin
      rob_uop_2_arch_dst <= _GEN_28934;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_2_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_2_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_2_dst_value <= _GEN_34056;
        end
      end else begin
        rob_uop_2_dst_value <= _GEN_34056;
      end
    end else begin
      rob_uop_2_dst_value <= _GEN_29638;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_2_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_2_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_2_src1_value <= _GEN_34120;
        end
      end else begin
        rob_uop_2_src1_value <= _GEN_34120;
      end
    end else begin
      rob_uop_2_src1_value <= _GEN_29702;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_2_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_2_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_2_alu_sel <= _GEN_34440;
        end
      end else begin
        rob_uop_2_alu_sel <= _GEN_34440;
      end
    end else begin
      rob_uop_2_alu_sel <= _GEN_30022;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_3_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_3_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_3_pc <= _GEN_32713;
        end
      end else begin
        rob_uop_3_pc <= _GEN_32713;
      end
    end else begin
      rob_uop_3_pc <= _GEN_28295;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_3_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_3_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_3_inst <= _GEN_32777;
        end
      end else begin
        rob_uop_3_inst <= _GEN_32777;
      end
    end else begin
      rob_uop_3_inst <= _GEN_28359;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_3_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_3_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_3_func_code <= _GEN_32841;
        end
      end else begin
        rob_uop_3_func_code <= _GEN_32841;
      end
    end else begin
      rob_uop_3_func_code <= _GEN_28423;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_3_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_3_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_3_phy_dst <= _GEN_33225;
        end
      end else begin
        rob_uop_3_phy_dst <= _GEN_33225;
      end
    end else begin
      rob_uop_3_phy_dst <= _GEN_28807;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_3_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_3_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_3_stale_dst <= _GEN_33289;
        end
      end else begin
        rob_uop_3_stale_dst <= _GEN_33289;
      end
    end else begin
      rob_uop_3_stale_dst <= _GEN_28871;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_3_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_3_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_3_arch_dst <= _GEN_33353;
        end
      end else begin
        rob_uop_3_arch_dst <= _GEN_33353;
      end
    end else begin
      rob_uop_3_arch_dst <= _GEN_28935;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_3_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_3_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_3_dst_value <= _GEN_34057;
        end
      end else begin
        rob_uop_3_dst_value <= _GEN_34057;
      end
    end else begin
      rob_uop_3_dst_value <= _GEN_29639;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_3_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_3_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_3_src1_value <= _GEN_34121;
        end
      end else begin
        rob_uop_3_src1_value <= _GEN_34121;
      end
    end else begin
      rob_uop_3_src1_value <= _GEN_29703;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_3_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_3_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_3_alu_sel <= _GEN_34441;
        end
      end else begin
        rob_uop_3_alu_sel <= _GEN_34441;
      end
    end else begin
      rob_uop_3_alu_sel <= _GEN_30023;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_4_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h4 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_4_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_4_pc <= _GEN_32714;
        end
      end else begin
        rob_uop_4_pc <= _GEN_32714;
      end
    end else begin
      rob_uop_4_pc <= _GEN_28296;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_4_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h4 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_4_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_4_inst <= _GEN_32778;
        end
      end else begin
        rob_uop_4_inst <= _GEN_32778;
      end
    end else begin
      rob_uop_4_inst <= _GEN_28360;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_4_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h4 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_4_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_4_func_code <= _GEN_32842;
        end
      end else begin
        rob_uop_4_func_code <= _GEN_32842;
      end
    end else begin
      rob_uop_4_func_code <= _GEN_28424;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_4_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h4 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_4_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_4_phy_dst <= _GEN_33226;
        end
      end else begin
        rob_uop_4_phy_dst <= _GEN_33226;
      end
    end else begin
      rob_uop_4_phy_dst <= _GEN_28808;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_4_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h4 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_4_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_4_stale_dst <= _GEN_33290;
        end
      end else begin
        rob_uop_4_stale_dst <= _GEN_33290;
      end
    end else begin
      rob_uop_4_stale_dst <= _GEN_28872;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_4_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h4 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_4_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_4_arch_dst <= _GEN_33354;
        end
      end else begin
        rob_uop_4_arch_dst <= _GEN_33354;
      end
    end else begin
      rob_uop_4_arch_dst <= _GEN_28936;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_4_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h4 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_4_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_4_dst_value <= _GEN_34058;
        end
      end else begin
        rob_uop_4_dst_value <= _GEN_34058;
      end
    end else begin
      rob_uop_4_dst_value <= _GEN_29640;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_4_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h4 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_4_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_4_src1_value <= _GEN_34122;
        end
      end else begin
        rob_uop_4_src1_value <= _GEN_34122;
      end
    end else begin
      rob_uop_4_src1_value <= _GEN_29704;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_4_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h4 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_4_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_4_alu_sel <= _GEN_34442;
        end
      end else begin
        rob_uop_4_alu_sel <= _GEN_34442;
      end
    end else begin
      rob_uop_4_alu_sel <= _GEN_30024;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_5_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h5 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_5_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_5_pc <= _GEN_32715;
        end
      end else begin
        rob_uop_5_pc <= _GEN_32715;
      end
    end else begin
      rob_uop_5_pc <= _GEN_28297;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_5_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h5 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_5_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_5_inst <= _GEN_32779;
        end
      end else begin
        rob_uop_5_inst <= _GEN_32779;
      end
    end else begin
      rob_uop_5_inst <= _GEN_28361;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_5_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h5 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_5_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_5_func_code <= _GEN_32843;
        end
      end else begin
        rob_uop_5_func_code <= _GEN_32843;
      end
    end else begin
      rob_uop_5_func_code <= _GEN_28425;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_5_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h5 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_5_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_5_phy_dst <= _GEN_33227;
        end
      end else begin
        rob_uop_5_phy_dst <= _GEN_33227;
      end
    end else begin
      rob_uop_5_phy_dst <= _GEN_28809;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_5_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h5 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_5_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_5_stale_dst <= _GEN_33291;
        end
      end else begin
        rob_uop_5_stale_dst <= _GEN_33291;
      end
    end else begin
      rob_uop_5_stale_dst <= _GEN_28873;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_5_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h5 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_5_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_5_arch_dst <= _GEN_33355;
        end
      end else begin
        rob_uop_5_arch_dst <= _GEN_33355;
      end
    end else begin
      rob_uop_5_arch_dst <= _GEN_28937;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_5_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h5 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_5_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_5_dst_value <= _GEN_34059;
        end
      end else begin
        rob_uop_5_dst_value <= _GEN_34059;
      end
    end else begin
      rob_uop_5_dst_value <= _GEN_29641;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_5_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h5 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_5_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_5_src1_value <= _GEN_34123;
        end
      end else begin
        rob_uop_5_src1_value <= _GEN_34123;
      end
    end else begin
      rob_uop_5_src1_value <= _GEN_29705;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_5_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h5 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_5_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_5_alu_sel <= _GEN_34443;
        end
      end else begin
        rob_uop_5_alu_sel <= _GEN_34443;
      end
    end else begin
      rob_uop_5_alu_sel <= _GEN_30025;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_6_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h6 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_6_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_6_pc <= _GEN_32716;
        end
      end else begin
        rob_uop_6_pc <= _GEN_32716;
      end
    end else begin
      rob_uop_6_pc <= _GEN_28298;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_6_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h6 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_6_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_6_inst <= _GEN_32780;
        end
      end else begin
        rob_uop_6_inst <= _GEN_32780;
      end
    end else begin
      rob_uop_6_inst <= _GEN_28362;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_6_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h6 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_6_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_6_func_code <= _GEN_32844;
        end
      end else begin
        rob_uop_6_func_code <= _GEN_32844;
      end
    end else begin
      rob_uop_6_func_code <= _GEN_28426;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_6_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h6 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_6_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_6_phy_dst <= _GEN_33228;
        end
      end else begin
        rob_uop_6_phy_dst <= _GEN_33228;
      end
    end else begin
      rob_uop_6_phy_dst <= _GEN_28810;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_6_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h6 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_6_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_6_stale_dst <= _GEN_33292;
        end
      end else begin
        rob_uop_6_stale_dst <= _GEN_33292;
      end
    end else begin
      rob_uop_6_stale_dst <= _GEN_28874;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_6_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h6 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_6_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_6_arch_dst <= _GEN_33356;
        end
      end else begin
        rob_uop_6_arch_dst <= _GEN_33356;
      end
    end else begin
      rob_uop_6_arch_dst <= _GEN_28938;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_6_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h6 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_6_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_6_dst_value <= _GEN_34060;
        end
      end else begin
        rob_uop_6_dst_value <= _GEN_34060;
      end
    end else begin
      rob_uop_6_dst_value <= _GEN_29642;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_6_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h6 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_6_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_6_src1_value <= _GEN_34124;
        end
      end else begin
        rob_uop_6_src1_value <= _GEN_34124;
      end
    end else begin
      rob_uop_6_src1_value <= _GEN_29706;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_6_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h6 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_6_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_6_alu_sel <= _GEN_34444;
        end
      end else begin
        rob_uop_6_alu_sel <= _GEN_34444;
      end
    end else begin
      rob_uop_6_alu_sel <= _GEN_30026;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_7_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h7 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_7_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_7_pc <= _GEN_32717;
        end
      end else begin
        rob_uop_7_pc <= _GEN_32717;
      end
    end else begin
      rob_uop_7_pc <= _GEN_28299;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_7_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h7 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_7_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_7_inst <= _GEN_32781;
        end
      end else begin
        rob_uop_7_inst <= _GEN_32781;
      end
    end else begin
      rob_uop_7_inst <= _GEN_28363;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_7_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h7 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_7_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_7_func_code <= _GEN_32845;
        end
      end else begin
        rob_uop_7_func_code <= _GEN_32845;
      end
    end else begin
      rob_uop_7_func_code <= _GEN_28427;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_7_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h7 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_7_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_7_phy_dst <= _GEN_33229;
        end
      end else begin
        rob_uop_7_phy_dst <= _GEN_33229;
      end
    end else begin
      rob_uop_7_phy_dst <= _GEN_28811;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_7_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h7 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_7_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_7_stale_dst <= _GEN_33293;
        end
      end else begin
        rob_uop_7_stale_dst <= _GEN_33293;
      end
    end else begin
      rob_uop_7_stale_dst <= _GEN_28875;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_7_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h7 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_7_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_7_arch_dst <= _GEN_33357;
        end
      end else begin
        rob_uop_7_arch_dst <= _GEN_33357;
      end
    end else begin
      rob_uop_7_arch_dst <= _GEN_28939;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_7_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h7 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_7_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_7_dst_value <= _GEN_34061;
        end
      end else begin
        rob_uop_7_dst_value <= _GEN_34061;
      end
    end else begin
      rob_uop_7_dst_value <= _GEN_29643;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_7_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h7 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_7_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_7_src1_value <= _GEN_34125;
        end
      end else begin
        rob_uop_7_src1_value <= _GEN_34125;
      end
    end else begin
      rob_uop_7_src1_value <= _GEN_29707;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_7_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h7 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_7_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_7_alu_sel <= _GEN_34445;
        end
      end else begin
        rob_uop_7_alu_sel <= _GEN_34445;
      end
    end else begin
      rob_uop_7_alu_sel <= _GEN_30027;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_8_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h8 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_8_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_8_pc <= _GEN_32718;
        end
      end else begin
        rob_uop_8_pc <= _GEN_32718;
      end
    end else begin
      rob_uop_8_pc <= _GEN_28300;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_8_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h8 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_8_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_8_inst <= _GEN_32782;
        end
      end else begin
        rob_uop_8_inst <= _GEN_32782;
      end
    end else begin
      rob_uop_8_inst <= _GEN_28364;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_8_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h8 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_8_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_8_func_code <= _GEN_32846;
        end
      end else begin
        rob_uop_8_func_code <= _GEN_32846;
      end
    end else begin
      rob_uop_8_func_code <= _GEN_28428;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_8_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h8 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_8_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_8_phy_dst <= _GEN_33230;
        end
      end else begin
        rob_uop_8_phy_dst <= _GEN_33230;
      end
    end else begin
      rob_uop_8_phy_dst <= _GEN_28812;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_8_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h8 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_8_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_8_stale_dst <= _GEN_33294;
        end
      end else begin
        rob_uop_8_stale_dst <= _GEN_33294;
      end
    end else begin
      rob_uop_8_stale_dst <= _GEN_28876;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_8_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h8 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_8_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_8_arch_dst <= _GEN_33358;
        end
      end else begin
        rob_uop_8_arch_dst <= _GEN_33358;
      end
    end else begin
      rob_uop_8_arch_dst <= _GEN_28940;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_8_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h8 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_8_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_8_dst_value <= _GEN_34062;
        end
      end else begin
        rob_uop_8_dst_value <= _GEN_34062;
      end
    end else begin
      rob_uop_8_dst_value <= _GEN_29644;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_8_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h8 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_8_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_8_src1_value <= _GEN_34126;
        end
      end else begin
        rob_uop_8_src1_value <= _GEN_34126;
      end
    end else begin
      rob_uop_8_src1_value <= _GEN_29708;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_8_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h8 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_8_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_8_alu_sel <= _GEN_34446;
        end
      end else begin
        rob_uop_8_alu_sel <= _GEN_34446;
      end
    end else begin
      rob_uop_8_alu_sel <= _GEN_30028;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_9_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h9 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_9_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_9_pc <= _GEN_32719;
        end
      end else begin
        rob_uop_9_pc <= _GEN_32719;
      end
    end else begin
      rob_uop_9_pc <= _GEN_28301;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_9_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h9 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_9_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_9_inst <= _GEN_32783;
        end
      end else begin
        rob_uop_9_inst <= _GEN_32783;
      end
    end else begin
      rob_uop_9_inst <= _GEN_28365;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_9_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h9 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_9_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_9_func_code <= _GEN_32847;
        end
      end else begin
        rob_uop_9_func_code <= _GEN_32847;
      end
    end else begin
      rob_uop_9_func_code <= _GEN_28429;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_9_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h9 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_9_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_9_phy_dst <= _GEN_33231;
        end
      end else begin
        rob_uop_9_phy_dst <= _GEN_33231;
      end
    end else begin
      rob_uop_9_phy_dst <= _GEN_28813;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_9_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h9 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_9_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_9_stale_dst <= _GEN_33295;
        end
      end else begin
        rob_uop_9_stale_dst <= _GEN_33295;
      end
    end else begin
      rob_uop_9_stale_dst <= _GEN_28877;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_9_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h9 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_9_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_9_arch_dst <= _GEN_33359;
        end
      end else begin
        rob_uop_9_arch_dst <= _GEN_33359;
      end
    end else begin
      rob_uop_9_arch_dst <= _GEN_28941;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_9_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h9 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_9_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_9_dst_value <= _GEN_34063;
        end
      end else begin
        rob_uop_9_dst_value <= _GEN_34063;
      end
    end else begin
      rob_uop_9_dst_value <= _GEN_29645;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_9_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h9 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_9_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_9_src1_value <= _GEN_34127;
        end
      end else begin
        rob_uop_9_src1_value <= _GEN_34127;
      end
    end else begin
      rob_uop_9_src1_value <= _GEN_29709;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_9_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h9 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_9_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_9_alu_sel <= _GEN_34447;
        end
      end else begin
        rob_uop_9_alu_sel <= _GEN_34447;
      end
    end else begin
      rob_uop_9_alu_sel <= _GEN_30029;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_10_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'ha == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_10_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_10_pc <= _GEN_32720;
        end
      end else begin
        rob_uop_10_pc <= _GEN_32720;
      end
    end else begin
      rob_uop_10_pc <= _GEN_28302;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_10_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'ha == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_10_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_10_inst <= _GEN_32784;
        end
      end else begin
        rob_uop_10_inst <= _GEN_32784;
      end
    end else begin
      rob_uop_10_inst <= _GEN_28366;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_10_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'ha == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_10_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_10_func_code <= _GEN_32848;
        end
      end else begin
        rob_uop_10_func_code <= _GEN_32848;
      end
    end else begin
      rob_uop_10_func_code <= _GEN_28430;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_10_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'ha == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_10_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_10_phy_dst <= _GEN_33232;
        end
      end else begin
        rob_uop_10_phy_dst <= _GEN_33232;
      end
    end else begin
      rob_uop_10_phy_dst <= _GEN_28814;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_10_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'ha == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_10_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_10_stale_dst <= _GEN_33296;
        end
      end else begin
        rob_uop_10_stale_dst <= _GEN_33296;
      end
    end else begin
      rob_uop_10_stale_dst <= _GEN_28878;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_10_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'ha == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_10_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_10_arch_dst <= _GEN_33360;
        end
      end else begin
        rob_uop_10_arch_dst <= _GEN_33360;
      end
    end else begin
      rob_uop_10_arch_dst <= _GEN_28942;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_10_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'ha == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_10_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_10_dst_value <= _GEN_34064;
        end
      end else begin
        rob_uop_10_dst_value <= _GEN_34064;
      end
    end else begin
      rob_uop_10_dst_value <= _GEN_29646;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_10_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'ha == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_10_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_10_src1_value <= _GEN_34128;
        end
      end else begin
        rob_uop_10_src1_value <= _GEN_34128;
      end
    end else begin
      rob_uop_10_src1_value <= _GEN_29710;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_10_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'ha == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_10_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_10_alu_sel <= _GEN_34448;
        end
      end else begin
        rob_uop_10_alu_sel <= _GEN_34448;
      end
    end else begin
      rob_uop_10_alu_sel <= _GEN_30030;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_11_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'hb == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_11_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_11_pc <= _GEN_32721;
        end
      end else begin
        rob_uop_11_pc <= _GEN_32721;
      end
    end else begin
      rob_uop_11_pc <= _GEN_28303;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_11_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'hb == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_11_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_11_inst <= _GEN_32785;
        end
      end else begin
        rob_uop_11_inst <= _GEN_32785;
      end
    end else begin
      rob_uop_11_inst <= _GEN_28367;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_11_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'hb == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_11_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_11_func_code <= _GEN_32849;
        end
      end else begin
        rob_uop_11_func_code <= _GEN_32849;
      end
    end else begin
      rob_uop_11_func_code <= _GEN_28431;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_11_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'hb == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_11_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_11_phy_dst <= _GEN_33233;
        end
      end else begin
        rob_uop_11_phy_dst <= _GEN_33233;
      end
    end else begin
      rob_uop_11_phy_dst <= _GEN_28815;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_11_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'hb == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_11_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_11_stale_dst <= _GEN_33297;
        end
      end else begin
        rob_uop_11_stale_dst <= _GEN_33297;
      end
    end else begin
      rob_uop_11_stale_dst <= _GEN_28879;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_11_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'hb == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_11_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_11_arch_dst <= _GEN_33361;
        end
      end else begin
        rob_uop_11_arch_dst <= _GEN_33361;
      end
    end else begin
      rob_uop_11_arch_dst <= _GEN_28943;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_11_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'hb == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_11_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_11_dst_value <= _GEN_34065;
        end
      end else begin
        rob_uop_11_dst_value <= _GEN_34065;
      end
    end else begin
      rob_uop_11_dst_value <= _GEN_29647;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_11_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'hb == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_11_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_11_src1_value <= _GEN_34129;
        end
      end else begin
        rob_uop_11_src1_value <= _GEN_34129;
      end
    end else begin
      rob_uop_11_src1_value <= _GEN_29711;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_11_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'hb == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_11_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_11_alu_sel <= _GEN_34449;
        end
      end else begin
        rob_uop_11_alu_sel <= _GEN_34449;
      end
    end else begin
      rob_uop_11_alu_sel <= _GEN_30031;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_12_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'hc == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_12_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_12_pc <= _GEN_32722;
        end
      end else begin
        rob_uop_12_pc <= _GEN_32722;
      end
    end else begin
      rob_uop_12_pc <= _GEN_28304;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_12_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'hc == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_12_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_12_inst <= _GEN_32786;
        end
      end else begin
        rob_uop_12_inst <= _GEN_32786;
      end
    end else begin
      rob_uop_12_inst <= _GEN_28368;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_12_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'hc == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_12_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_12_func_code <= _GEN_32850;
        end
      end else begin
        rob_uop_12_func_code <= _GEN_32850;
      end
    end else begin
      rob_uop_12_func_code <= _GEN_28432;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_12_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'hc == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_12_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_12_phy_dst <= _GEN_33234;
        end
      end else begin
        rob_uop_12_phy_dst <= _GEN_33234;
      end
    end else begin
      rob_uop_12_phy_dst <= _GEN_28816;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_12_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'hc == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_12_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_12_stale_dst <= _GEN_33298;
        end
      end else begin
        rob_uop_12_stale_dst <= _GEN_33298;
      end
    end else begin
      rob_uop_12_stale_dst <= _GEN_28880;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_12_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'hc == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_12_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_12_arch_dst <= _GEN_33362;
        end
      end else begin
        rob_uop_12_arch_dst <= _GEN_33362;
      end
    end else begin
      rob_uop_12_arch_dst <= _GEN_28944;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_12_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'hc == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_12_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_12_dst_value <= _GEN_34066;
        end
      end else begin
        rob_uop_12_dst_value <= _GEN_34066;
      end
    end else begin
      rob_uop_12_dst_value <= _GEN_29648;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_12_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'hc == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_12_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_12_src1_value <= _GEN_34130;
        end
      end else begin
        rob_uop_12_src1_value <= _GEN_34130;
      end
    end else begin
      rob_uop_12_src1_value <= _GEN_29712;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_12_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'hc == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_12_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_12_alu_sel <= _GEN_34450;
        end
      end else begin
        rob_uop_12_alu_sel <= _GEN_34450;
      end
    end else begin
      rob_uop_12_alu_sel <= _GEN_30032;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_13_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'hd == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_13_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_13_pc <= _GEN_32723;
        end
      end else begin
        rob_uop_13_pc <= _GEN_32723;
      end
    end else begin
      rob_uop_13_pc <= _GEN_28305;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_13_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'hd == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_13_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_13_inst <= _GEN_32787;
        end
      end else begin
        rob_uop_13_inst <= _GEN_32787;
      end
    end else begin
      rob_uop_13_inst <= _GEN_28369;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_13_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'hd == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_13_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_13_func_code <= _GEN_32851;
        end
      end else begin
        rob_uop_13_func_code <= _GEN_32851;
      end
    end else begin
      rob_uop_13_func_code <= _GEN_28433;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_13_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'hd == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_13_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_13_phy_dst <= _GEN_33235;
        end
      end else begin
        rob_uop_13_phy_dst <= _GEN_33235;
      end
    end else begin
      rob_uop_13_phy_dst <= _GEN_28817;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_13_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'hd == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_13_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_13_stale_dst <= _GEN_33299;
        end
      end else begin
        rob_uop_13_stale_dst <= _GEN_33299;
      end
    end else begin
      rob_uop_13_stale_dst <= _GEN_28881;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_13_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'hd == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_13_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_13_arch_dst <= _GEN_33363;
        end
      end else begin
        rob_uop_13_arch_dst <= _GEN_33363;
      end
    end else begin
      rob_uop_13_arch_dst <= _GEN_28945;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_13_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'hd == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_13_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_13_dst_value <= _GEN_34067;
        end
      end else begin
        rob_uop_13_dst_value <= _GEN_34067;
      end
    end else begin
      rob_uop_13_dst_value <= _GEN_29649;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_13_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'hd == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_13_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_13_src1_value <= _GEN_34131;
        end
      end else begin
        rob_uop_13_src1_value <= _GEN_34131;
      end
    end else begin
      rob_uop_13_src1_value <= _GEN_29713;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_13_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'hd == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_13_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_13_alu_sel <= _GEN_34451;
        end
      end else begin
        rob_uop_13_alu_sel <= _GEN_34451;
      end
    end else begin
      rob_uop_13_alu_sel <= _GEN_30033;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_14_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'he == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_14_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_14_pc <= _GEN_32724;
        end
      end else begin
        rob_uop_14_pc <= _GEN_32724;
      end
    end else begin
      rob_uop_14_pc <= _GEN_28306;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_14_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'he == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_14_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_14_inst <= _GEN_32788;
        end
      end else begin
        rob_uop_14_inst <= _GEN_32788;
      end
    end else begin
      rob_uop_14_inst <= _GEN_28370;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_14_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'he == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_14_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_14_func_code <= _GEN_32852;
        end
      end else begin
        rob_uop_14_func_code <= _GEN_32852;
      end
    end else begin
      rob_uop_14_func_code <= _GEN_28434;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_14_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'he == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_14_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_14_phy_dst <= _GEN_33236;
        end
      end else begin
        rob_uop_14_phy_dst <= _GEN_33236;
      end
    end else begin
      rob_uop_14_phy_dst <= _GEN_28818;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_14_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'he == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_14_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_14_stale_dst <= _GEN_33300;
        end
      end else begin
        rob_uop_14_stale_dst <= _GEN_33300;
      end
    end else begin
      rob_uop_14_stale_dst <= _GEN_28882;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_14_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'he == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_14_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_14_arch_dst <= _GEN_33364;
        end
      end else begin
        rob_uop_14_arch_dst <= _GEN_33364;
      end
    end else begin
      rob_uop_14_arch_dst <= _GEN_28946;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_14_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'he == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_14_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_14_dst_value <= _GEN_34068;
        end
      end else begin
        rob_uop_14_dst_value <= _GEN_34068;
      end
    end else begin
      rob_uop_14_dst_value <= _GEN_29650;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_14_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'he == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_14_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_14_src1_value <= _GEN_34132;
        end
      end else begin
        rob_uop_14_src1_value <= _GEN_34132;
      end
    end else begin
      rob_uop_14_src1_value <= _GEN_29714;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_14_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'he == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_14_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_14_alu_sel <= _GEN_34452;
        end
      end else begin
        rob_uop_14_alu_sel <= _GEN_34452;
      end
    end else begin
      rob_uop_14_alu_sel <= _GEN_30034;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_15_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'hf == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_15_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_15_pc <= _GEN_32725;
        end
      end else begin
        rob_uop_15_pc <= _GEN_32725;
      end
    end else begin
      rob_uop_15_pc <= _GEN_28307;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_15_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'hf == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_15_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_15_inst <= _GEN_32789;
        end
      end else begin
        rob_uop_15_inst <= _GEN_32789;
      end
    end else begin
      rob_uop_15_inst <= _GEN_28371;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_15_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'hf == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_15_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_15_func_code <= _GEN_32853;
        end
      end else begin
        rob_uop_15_func_code <= _GEN_32853;
      end
    end else begin
      rob_uop_15_func_code <= _GEN_28435;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_15_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'hf == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_15_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_15_phy_dst <= _GEN_33237;
        end
      end else begin
        rob_uop_15_phy_dst <= _GEN_33237;
      end
    end else begin
      rob_uop_15_phy_dst <= _GEN_28819;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_15_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'hf == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_15_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_15_stale_dst <= _GEN_33301;
        end
      end else begin
        rob_uop_15_stale_dst <= _GEN_33301;
      end
    end else begin
      rob_uop_15_stale_dst <= _GEN_28883;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_15_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'hf == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_15_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_15_arch_dst <= _GEN_33365;
        end
      end else begin
        rob_uop_15_arch_dst <= _GEN_33365;
      end
    end else begin
      rob_uop_15_arch_dst <= _GEN_28947;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_15_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'hf == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_15_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_15_dst_value <= _GEN_34069;
        end
      end else begin
        rob_uop_15_dst_value <= _GEN_34069;
      end
    end else begin
      rob_uop_15_dst_value <= _GEN_29651;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_15_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'hf == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_15_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_15_src1_value <= _GEN_34133;
        end
      end else begin
        rob_uop_15_src1_value <= _GEN_34133;
      end
    end else begin
      rob_uop_15_src1_value <= _GEN_29715;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_15_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'hf == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_15_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_15_alu_sel <= _GEN_34453;
        end
      end else begin
        rob_uop_15_alu_sel <= _GEN_34453;
      end
    end else begin
      rob_uop_15_alu_sel <= _GEN_30035;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_16_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h10 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_16_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_16_pc <= _GEN_32726;
        end
      end else begin
        rob_uop_16_pc <= _GEN_32726;
      end
    end else begin
      rob_uop_16_pc <= _GEN_28308;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_16_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h10 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_16_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_16_inst <= _GEN_32790;
        end
      end else begin
        rob_uop_16_inst <= _GEN_32790;
      end
    end else begin
      rob_uop_16_inst <= _GEN_28372;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_16_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h10 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_16_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_16_func_code <= _GEN_32854;
        end
      end else begin
        rob_uop_16_func_code <= _GEN_32854;
      end
    end else begin
      rob_uop_16_func_code <= _GEN_28436;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_16_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h10 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_16_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_16_phy_dst <= _GEN_33238;
        end
      end else begin
        rob_uop_16_phy_dst <= _GEN_33238;
      end
    end else begin
      rob_uop_16_phy_dst <= _GEN_28820;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_16_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h10 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_16_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_16_stale_dst <= _GEN_33302;
        end
      end else begin
        rob_uop_16_stale_dst <= _GEN_33302;
      end
    end else begin
      rob_uop_16_stale_dst <= _GEN_28884;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_16_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h10 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_16_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_16_arch_dst <= _GEN_33366;
        end
      end else begin
        rob_uop_16_arch_dst <= _GEN_33366;
      end
    end else begin
      rob_uop_16_arch_dst <= _GEN_28948;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_16_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h10 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_16_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_16_dst_value <= _GEN_34070;
        end
      end else begin
        rob_uop_16_dst_value <= _GEN_34070;
      end
    end else begin
      rob_uop_16_dst_value <= _GEN_29652;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_16_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h10 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_16_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_16_src1_value <= _GEN_34134;
        end
      end else begin
        rob_uop_16_src1_value <= _GEN_34134;
      end
    end else begin
      rob_uop_16_src1_value <= _GEN_29716;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_16_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h10 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_16_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_16_alu_sel <= _GEN_34454;
        end
      end else begin
        rob_uop_16_alu_sel <= _GEN_34454;
      end
    end else begin
      rob_uop_16_alu_sel <= _GEN_30036;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_17_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h11 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_17_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_17_pc <= _GEN_32727;
        end
      end else begin
        rob_uop_17_pc <= _GEN_32727;
      end
    end else begin
      rob_uop_17_pc <= _GEN_28309;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_17_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h11 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_17_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_17_inst <= _GEN_32791;
        end
      end else begin
        rob_uop_17_inst <= _GEN_32791;
      end
    end else begin
      rob_uop_17_inst <= _GEN_28373;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_17_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h11 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_17_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_17_func_code <= _GEN_32855;
        end
      end else begin
        rob_uop_17_func_code <= _GEN_32855;
      end
    end else begin
      rob_uop_17_func_code <= _GEN_28437;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_17_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h11 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_17_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_17_phy_dst <= _GEN_33239;
        end
      end else begin
        rob_uop_17_phy_dst <= _GEN_33239;
      end
    end else begin
      rob_uop_17_phy_dst <= _GEN_28821;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_17_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h11 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_17_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_17_stale_dst <= _GEN_33303;
        end
      end else begin
        rob_uop_17_stale_dst <= _GEN_33303;
      end
    end else begin
      rob_uop_17_stale_dst <= _GEN_28885;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_17_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h11 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_17_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_17_arch_dst <= _GEN_33367;
        end
      end else begin
        rob_uop_17_arch_dst <= _GEN_33367;
      end
    end else begin
      rob_uop_17_arch_dst <= _GEN_28949;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_17_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h11 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_17_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_17_dst_value <= _GEN_34071;
        end
      end else begin
        rob_uop_17_dst_value <= _GEN_34071;
      end
    end else begin
      rob_uop_17_dst_value <= _GEN_29653;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_17_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h11 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_17_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_17_src1_value <= _GEN_34135;
        end
      end else begin
        rob_uop_17_src1_value <= _GEN_34135;
      end
    end else begin
      rob_uop_17_src1_value <= _GEN_29717;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_17_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h11 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_17_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_17_alu_sel <= _GEN_34455;
        end
      end else begin
        rob_uop_17_alu_sel <= _GEN_34455;
      end
    end else begin
      rob_uop_17_alu_sel <= _GEN_30037;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_18_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h12 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_18_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_18_pc <= _GEN_32728;
        end
      end else begin
        rob_uop_18_pc <= _GEN_32728;
      end
    end else begin
      rob_uop_18_pc <= _GEN_28310;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_18_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h12 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_18_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_18_inst <= _GEN_32792;
        end
      end else begin
        rob_uop_18_inst <= _GEN_32792;
      end
    end else begin
      rob_uop_18_inst <= _GEN_28374;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_18_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h12 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_18_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_18_func_code <= _GEN_32856;
        end
      end else begin
        rob_uop_18_func_code <= _GEN_32856;
      end
    end else begin
      rob_uop_18_func_code <= _GEN_28438;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_18_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h12 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_18_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_18_phy_dst <= _GEN_33240;
        end
      end else begin
        rob_uop_18_phy_dst <= _GEN_33240;
      end
    end else begin
      rob_uop_18_phy_dst <= _GEN_28822;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_18_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h12 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_18_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_18_stale_dst <= _GEN_33304;
        end
      end else begin
        rob_uop_18_stale_dst <= _GEN_33304;
      end
    end else begin
      rob_uop_18_stale_dst <= _GEN_28886;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_18_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h12 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_18_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_18_arch_dst <= _GEN_33368;
        end
      end else begin
        rob_uop_18_arch_dst <= _GEN_33368;
      end
    end else begin
      rob_uop_18_arch_dst <= _GEN_28950;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_18_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h12 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_18_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_18_dst_value <= _GEN_34072;
        end
      end else begin
        rob_uop_18_dst_value <= _GEN_34072;
      end
    end else begin
      rob_uop_18_dst_value <= _GEN_29654;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_18_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h12 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_18_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_18_src1_value <= _GEN_34136;
        end
      end else begin
        rob_uop_18_src1_value <= _GEN_34136;
      end
    end else begin
      rob_uop_18_src1_value <= _GEN_29718;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_18_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h12 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_18_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_18_alu_sel <= _GEN_34456;
        end
      end else begin
        rob_uop_18_alu_sel <= _GEN_34456;
      end
    end else begin
      rob_uop_18_alu_sel <= _GEN_30038;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_19_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h13 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_19_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_19_pc <= _GEN_32729;
        end
      end else begin
        rob_uop_19_pc <= _GEN_32729;
      end
    end else begin
      rob_uop_19_pc <= _GEN_28311;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_19_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h13 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_19_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_19_inst <= _GEN_32793;
        end
      end else begin
        rob_uop_19_inst <= _GEN_32793;
      end
    end else begin
      rob_uop_19_inst <= _GEN_28375;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_19_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h13 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_19_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_19_func_code <= _GEN_32857;
        end
      end else begin
        rob_uop_19_func_code <= _GEN_32857;
      end
    end else begin
      rob_uop_19_func_code <= _GEN_28439;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_19_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h13 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_19_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_19_phy_dst <= _GEN_33241;
        end
      end else begin
        rob_uop_19_phy_dst <= _GEN_33241;
      end
    end else begin
      rob_uop_19_phy_dst <= _GEN_28823;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_19_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h13 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_19_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_19_stale_dst <= _GEN_33305;
        end
      end else begin
        rob_uop_19_stale_dst <= _GEN_33305;
      end
    end else begin
      rob_uop_19_stale_dst <= _GEN_28887;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_19_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h13 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_19_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_19_arch_dst <= _GEN_33369;
        end
      end else begin
        rob_uop_19_arch_dst <= _GEN_33369;
      end
    end else begin
      rob_uop_19_arch_dst <= _GEN_28951;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_19_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h13 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_19_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_19_dst_value <= _GEN_34073;
        end
      end else begin
        rob_uop_19_dst_value <= _GEN_34073;
      end
    end else begin
      rob_uop_19_dst_value <= _GEN_29655;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_19_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h13 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_19_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_19_src1_value <= _GEN_34137;
        end
      end else begin
        rob_uop_19_src1_value <= _GEN_34137;
      end
    end else begin
      rob_uop_19_src1_value <= _GEN_29719;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_19_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h13 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_19_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_19_alu_sel <= _GEN_34457;
        end
      end else begin
        rob_uop_19_alu_sel <= _GEN_34457;
      end
    end else begin
      rob_uop_19_alu_sel <= _GEN_30039;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_20_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h14 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_20_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_20_pc <= _GEN_32730;
        end
      end else begin
        rob_uop_20_pc <= _GEN_32730;
      end
    end else begin
      rob_uop_20_pc <= _GEN_28312;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_20_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h14 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_20_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_20_inst <= _GEN_32794;
        end
      end else begin
        rob_uop_20_inst <= _GEN_32794;
      end
    end else begin
      rob_uop_20_inst <= _GEN_28376;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_20_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h14 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_20_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_20_func_code <= _GEN_32858;
        end
      end else begin
        rob_uop_20_func_code <= _GEN_32858;
      end
    end else begin
      rob_uop_20_func_code <= _GEN_28440;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_20_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h14 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_20_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_20_phy_dst <= _GEN_33242;
        end
      end else begin
        rob_uop_20_phy_dst <= _GEN_33242;
      end
    end else begin
      rob_uop_20_phy_dst <= _GEN_28824;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_20_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h14 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_20_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_20_stale_dst <= _GEN_33306;
        end
      end else begin
        rob_uop_20_stale_dst <= _GEN_33306;
      end
    end else begin
      rob_uop_20_stale_dst <= _GEN_28888;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_20_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h14 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_20_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_20_arch_dst <= _GEN_33370;
        end
      end else begin
        rob_uop_20_arch_dst <= _GEN_33370;
      end
    end else begin
      rob_uop_20_arch_dst <= _GEN_28952;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_20_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h14 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_20_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_20_dst_value <= _GEN_34074;
        end
      end else begin
        rob_uop_20_dst_value <= _GEN_34074;
      end
    end else begin
      rob_uop_20_dst_value <= _GEN_29656;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_20_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h14 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_20_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_20_src1_value <= _GEN_34138;
        end
      end else begin
        rob_uop_20_src1_value <= _GEN_34138;
      end
    end else begin
      rob_uop_20_src1_value <= _GEN_29720;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_20_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h14 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_20_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_20_alu_sel <= _GEN_34458;
        end
      end else begin
        rob_uop_20_alu_sel <= _GEN_34458;
      end
    end else begin
      rob_uop_20_alu_sel <= _GEN_30040;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_21_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h15 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_21_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_21_pc <= _GEN_32731;
        end
      end else begin
        rob_uop_21_pc <= _GEN_32731;
      end
    end else begin
      rob_uop_21_pc <= _GEN_28313;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_21_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h15 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_21_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_21_inst <= _GEN_32795;
        end
      end else begin
        rob_uop_21_inst <= _GEN_32795;
      end
    end else begin
      rob_uop_21_inst <= _GEN_28377;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_21_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h15 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_21_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_21_func_code <= _GEN_32859;
        end
      end else begin
        rob_uop_21_func_code <= _GEN_32859;
      end
    end else begin
      rob_uop_21_func_code <= _GEN_28441;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_21_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h15 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_21_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_21_phy_dst <= _GEN_33243;
        end
      end else begin
        rob_uop_21_phy_dst <= _GEN_33243;
      end
    end else begin
      rob_uop_21_phy_dst <= _GEN_28825;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_21_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h15 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_21_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_21_stale_dst <= _GEN_33307;
        end
      end else begin
        rob_uop_21_stale_dst <= _GEN_33307;
      end
    end else begin
      rob_uop_21_stale_dst <= _GEN_28889;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_21_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h15 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_21_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_21_arch_dst <= _GEN_33371;
        end
      end else begin
        rob_uop_21_arch_dst <= _GEN_33371;
      end
    end else begin
      rob_uop_21_arch_dst <= _GEN_28953;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_21_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h15 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_21_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_21_dst_value <= _GEN_34075;
        end
      end else begin
        rob_uop_21_dst_value <= _GEN_34075;
      end
    end else begin
      rob_uop_21_dst_value <= _GEN_29657;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_21_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h15 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_21_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_21_src1_value <= _GEN_34139;
        end
      end else begin
        rob_uop_21_src1_value <= _GEN_34139;
      end
    end else begin
      rob_uop_21_src1_value <= _GEN_29721;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_21_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h15 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_21_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_21_alu_sel <= _GEN_34459;
        end
      end else begin
        rob_uop_21_alu_sel <= _GEN_34459;
      end
    end else begin
      rob_uop_21_alu_sel <= _GEN_30041;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_22_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h16 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_22_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_22_pc <= _GEN_32732;
        end
      end else begin
        rob_uop_22_pc <= _GEN_32732;
      end
    end else begin
      rob_uop_22_pc <= _GEN_28314;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_22_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h16 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_22_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_22_inst <= _GEN_32796;
        end
      end else begin
        rob_uop_22_inst <= _GEN_32796;
      end
    end else begin
      rob_uop_22_inst <= _GEN_28378;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_22_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h16 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_22_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_22_func_code <= _GEN_32860;
        end
      end else begin
        rob_uop_22_func_code <= _GEN_32860;
      end
    end else begin
      rob_uop_22_func_code <= _GEN_28442;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_22_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h16 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_22_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_22_phy_dst <= _GEN_33244;
        end
      end else begin
        rob_uop_22_phy_dst <= _GEN_33244;
      end
    end else begin
      rob_uop_22_phy_dst <= _GEN_28826;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_22_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h16 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_22_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_22_stale_dst <= _GEN_33308;
        end
      end else begin
        rob_uop_22_stale_dst <= _GEN_33308;
      end
    end else begin
      rob_uop_22_stale_dst <= _GEN_28890;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_22_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h16 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_22_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_22_arch_dst <= _GEN_33372;
        end
      end else begin
        rob_uop_22_arch_dst <= _GEN_33372;
      end
    end else begin
      rob_uop_22_arch_dst <= _GEN_28954;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_22_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h16 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_22_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_22_dst_value <= _GEN_34076;
        end
      end else begin
        rob_uop_22_dst_value <= _GEN_34076;
      end
    end else begin
      rob_uop_22_dst_value <= _GEN_29658;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_22_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h16 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_22_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_22_src1_value <= _GEN_34140;
        end
      end else begin
        rob_uop_22_src1_value <= _GEN_34140;
      end
    end else begin
      rob_uop_22_src1_value <= _GEN_29722;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_22_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h16 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_22_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_22_alu_sel <= _GEN_34460;
        end
      end else begin
        rob_uop_22_alu_sel <= _GEN_34460;
      end
    end else begin
      rob_uop_22_alu_sel <= _GEN_30042;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_23_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h17 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_23_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_23_pc <= _GEN_32733;
        end
      end else begin
        rob_uop_23_pc <= _GEN_32733;
      end
    end else begin
      rob_uop_23_pc <= _GEN_28315;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_23_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h17 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_23_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_23_inst <= _GEN_32797;
        end
      end else begin
        rob_uop_23_inst <= _GEN_32797;
      end
    end else begin
      rob_uop_23_inst <= _GEN_28379;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_23_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h17 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_23_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_23_func_code <= _GEN_32861;
        end
      end else begin
        rob_uop_23_func_code <= _GEN_32861;
      end
    end else begin
      rob_uop_23_func_code <= _GEN_28443;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_23_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h17 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_23_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_23_phy_dst <= _GEN_33245;
        end
      end else begin
        rob_uop_23_phy_dst <= _GEN_33245;
      end
    end else begin
      rob_uop_23_phy_dst <= _GEN_28827;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_23_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h17 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_23_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_23_stale_dst <= _GEN_33309;
        end
      end else begin
        rob_uop_23_stale_dst <= _GEN_33309;
      end
    end else begin
      rob_uop_23_stale_dst <= _GEN_28891;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_23_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h17 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_23_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_23_arch_dst <= _GEN_33373;
        end
      end else begin
        rob_uop_23_arch_dst <= _GEN_33373;
      end
    end else begin
      rob_uop_23_arch_dst <= _GEN_28955;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_23_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h17 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_23_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_23_dst_value <= _GEN_34077;
        end
      end else begin
        rob_uop_23_dst_value <= _GEN_34077;
      end
    end else begin
      rob_uop_23_dst_value <= _GEN_29659;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_23_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h17 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_23_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_23_src1_value <= _GEN_34141;
        end
      end else begin
        rob_uop_23_src1_value <= _GEN_34141;
      end
    end else begin
      rob_uop_23_src1_value <= _GEN_29723;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_23_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h17 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_23_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_23_alu_sel <= _GEN_34461;
        end
      end else begin
        rob_uop_23_alu_sel <= _GEN_34461;
      end
    end else begin
      rob_uop_23_alu_sel <= _GEN_30043;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_24_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h18 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_24_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_24_pc <= _GEN_32734;
        end
      end else begin
        rob_uop_24_pc <= _GEN_32734;
      end
    end else begin
      rob_uop_24_pc <= _GEN_28316;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_24_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h18 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_24_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_24_inst <= _GEN_32798;
        end
      end else begin
        rob_uop_24_inst <= _GEN_32798;
      end
    end else begin
      rob_uop_24_inst <= _GEN_28380;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_24_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h18 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_24_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_24_func_code <= _GEN_32862;
        end
      end else begin
        rob_uop_24_func_code <= _GEN_32862;
      end
    end else begin
      rob_uop_24_func_code <= _GEN_28444;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_24_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h18 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_24_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_24_phy_dst <= _GEN_33246;
        end
      end else begin
        rob_uop_24_phy_dst <= _GEN_33246;
      end
    end else begin
      rob_uop_24_phy_dst <= _GEN_28828;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_24_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h18 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_24_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_24_stale_dst <= _GEN_33310;
        end
      end else begin
        rob_uop_24_stale_dst <= _GEN_33310;
      end
    end else begin
      rob_uop_24_stale_dst <= _GEN_28892;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_24_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h18 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_24_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_24_arch_dst <= _GEN_33374;
        end
      end else begin
        rob_uop_24_arch_dst <= _GEN_33374;
      end
    end else begin
      rob_uop_24_arch_dst <= _GEN_28956;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_24_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h18 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_24_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_24_dst_value <= _GEN_34078;
        end
      end else begin
        rob_uop_24_dst_value <= _GEN_34078;
      end
    end else begin
      rob_uop_24_dst_value <= _GEN_29660;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_24_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h18 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_24_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_24_src1_value <= _GEN_34142;
        end
      end else begin
        rob_uop_24_src1_value <= _GEN_34142;
      end
    end else begin
      rob_uop_24_src1_value <= _GEN_29724;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_24_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h18 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_24_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_24_alu_sel <= _GEN_34462;
        end
      end else begin
        rob_uop_24_alu_sel <= _GEN_34462;
      end
    end else begin
      rob_uop_24_alu_sel <= _GEN_30044;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_25_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h19 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_25_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_25_pc <= _GEN_32735;
        end
      end else begin
        rob_uop_25_pc <= _GEN_32735;
      end
    end else begin
      rob_uop_25_pc <= _GEN_28317;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_25_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h19 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_25_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_25_inst <= _GEN_32799;
        end
      end else begin
        rob_uop_25_inst <= _GEN_32799;
      end
    end else begin
      rob_uop_25_inst <= _GEN_28381;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_25_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h19 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_25_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_25_func_code <= _GEN_32863;
        end
      end else begin
        rob_uop_25_func_code <= _GEN_32863;
      end
    end else begin
      rob_uop_25_func_code <= _GEN_28445;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_25_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h19 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_25_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_25_phy_dst <= _GEN_33247;
        end
      end else begin
        rob_uop_25_phy_dst <= _GEN_33247;
      end
    end else begin
      rob_uop_25_phy_dst <= _GEN_28829;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_25_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h19 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_25_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_25_stale_dst <= _GEN_33311;
        end
      end else begin
        rob_uop_25_stale_dst <= _GEN_33311;
      end
    end else begin
      rob_uop_25_stale_dst <= _GEN_28893;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_25_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h19 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_25_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_25_arch_dst <= _GEN_33375;
        end
      end else begin
        rob_uop_25_arch_dst <= _GEN_33375;
      end
    end else begin
      rob_uop_25_arch_dst <= _GEN_28957;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_25_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h19 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_25_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_25_dst_value <= _GEN_34079;
        end
      end else begin
        rob_uop_25_dst_value <= _GEN_34079;
      end
    end else begin
      rob_uop_25_dst_value <= _GEN_29661;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_25_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h19 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_25_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_25_src1_value <= _GEN_34143;
        end
      end else begin
        rob_uop_25_src1_value <= _GEN_34143;
      end
    end else begin
      rob_uop_25_src1_value <= _GEN_29725;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_25_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h19 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_25_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_25_alu_sel <= _GEN_34463;
        end
      end else begin
        rob_uop_25_alu_sel <= _GEN_34463;
      end
    end else begin
      rob_uop_25_alu_sel <= _GEN_30045;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_26_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1a == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_26_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_26_pc <= _GEN_32736;
        end
      end else begin
        rob_uop_26_pc <= _GEN_32736;
      end
    end else begin
      rob_uop_26_pc <= _GEN_28318;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_26_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1a == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_26_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_26_inst <= _GEN_32800;
        end
      end else begin
        rob_uop_26_inst <= _GEN_32800;
      end
    end else begin
      rob_uop_26_inst <= _GEN_28382;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_26_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1a == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_26_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_26_func_code <= _GEN_32864;
        end
      end else begin
        rob_uop_26_func_code <= _GEN_32864;
      end
    end else begin
      rob_uop_26_func_code <= _GEN_28446;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_26_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1a == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_26_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_26_phy_dst <= _GEN_33248;
        end
      end else begin
        rob_uop_26_phy_dst <= _GEN_33248;
      end
    end else begin
      rob_uop_26_phy_dst <= _GEN_28830;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_26_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1a == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_26_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_26_stale_dst <= _GEN_33312;
        end
      end else begin
        rob_uop_26_stale_dst <= _GEN_33312;
      end
    end else begin
      rob_uop_26_stale_dst <= _GEN_28894;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_26_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1a == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_26_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_26_arch_dst <= _GEN_33376;
        end
      end else begin
        rob_uop_26_arch_dst <= _GEN_33376;
      end
    end else begin
      rob_uop_26_arch_dst <= _GEN_28958;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_26_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1a == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_26_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_26_dst_value <= _GEN_34080;
        end
      end else begin
        rob_uop_26_dst_value <= _GEN_34080;
      end
    end else begin
      rob_uop_26_dst_value <= _GEN_29662;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_26_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1a == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_26_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_26_src1_value <= _GEN_34144;
        end
      end else begin
        rob_uop_26_src1_value <= _GEN_34144;
      end
    end else begin
      rob_uop_26_src1_value <= _GEN_29726;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_26_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1a == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_26_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_26_alu_sel <= _GEN_34464;
        end
      end else begin
        rob_uop_26_alu_sel <= _GEN_34464;
      end
    end else begin
      rob_uop_26_alu_sel <= _GEN_30046;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_27_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1b == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_27_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_27_pc <= _GEN_32737;
        end
      end else begin
        rob_uop_27_pc <= _GEN_32737;
      end
    end else begin
      rob_uop_27_pc <= _GEN_28319;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_27_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1b == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_27_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_27_inst <= _GEN_32801;
        end
      end else begin
        rob_uop_27_inst <= _GEN_32801;
      end
    end else begin
      rob_uop_27_inst <= _GEN_28383;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_27_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1b == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_27_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_27_func_code <= _GEN_32865;
        end
      end else begin
        rob_uop_27_func_code <= _GEN_32865;
      end
    end else begin
      rob_uop_27_func_code <= _GEN_28447;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_27_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1b == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_27_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_27_phy_dst <= _GEN_33249;
        end
      end else begin
        rob_uop_27_phy_dst <= _GEN_33249;
      end
    end else begin
      rob_uop_27_phy_dst <= _GEN_28831;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_27_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1b == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_27_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_27_stale_dst <= _GEN_33313;
        end
      end else begin
        rob_uop_27_stale_dst <= _GEN_33313;
      end
    end else begin
      rob_uop_27_stale_dst <= _GEN_28895;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_27_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1b == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_27_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_27_arch_dst <= _GEN_33377;
        end
      end else begin
        rob_uop_27_arch_dst <= _GEN_33377;
      end
    end else begin
      rob_uop_27_arch_dst <= _GEN_28959;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_27_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1b == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_27_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_27_dst_value <= _GEN_34081;
        end
      end else begin
        rob_uop_27_dst_value <= _GEN_34081;
      end
    end else begin
      rob_uop_27_dst_value <= _GEN_29663;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_27_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1b == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_27_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_27_src1_value <= _GEN_34145;
        end
      end else begin
        rob_uop_27_src1_value <= _GEN_34145;
      end
    end else begin
      rob_uop_27_src1_value <= _GEN_29727;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_27_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1b == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_27_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_27_alu_sel <= _GEN_34465;
        end
      end else begin
        rob_uop_27_alu_sel <= _GEN_34465;
      end
    end else begin
      rob_uop_27_alu_sel <= _GEN_30047;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_28_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1c == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_28_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_28_pc <= _GEN_32738;
        end
      end else begin
        rob_uop_28_pc <= _GEN_32738;
      end
    end else begin
      rob_uop_28_pc <= _GEN_28320;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_28_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1c == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_28_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_28_inst <= _GEN_32802;
        end
      end else begin
        rob_uop_28_inst <= _GEN_32802;
      end
    end else begin
      rob_uop_28_inst <= _GEN_28384;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_28_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1c == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_28_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_28_func_code <= _GEN_32866;
        end
      end else begin
        rob_uop_28_func_code <= _GEN_32866;
      end
    end else begin
      rob_uop_28_func_code <= _GEN_28448;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_28_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1c == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_28_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_28_phy_dst <= _GEN_33250;
        end
      end else begin
        rob_uop_28_phy_dst <= _GEN_33250;
      end
    end else begin
      rob_uop_28_phy_dst <= _GEN_28832;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_28_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1c == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_28_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_28_stale_dst <= _GEN_33314;
        end
      end else begin
        rob_uop_28_stale_dst <= _GEN_33314;
      end
    end else begin
      rob_uop_28_stale_dst <= _GEN_28896;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_28_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1c == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_28_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_28_arch_dst <= _GEN_33378;
        end
      end else begin
        rob_uop_28_arch_dst <= _GEN_33378;
      end
    end else begin
      rob_uop_28_arch_dst <= _GEN_28960;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_28_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1c == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_28_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_28_dst_value <= _GEN_34082;
        end
      end else begin
        rob_uop_28_dst_value <= _GEN_34082;
      end
    end else begin
      rob_uop_28_dst_value <= _GEN_29664;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_28_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1c == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_28_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_28_src1_value <= _GEN_34146;
        end
      end else begin
        rob_uop_28_src1_value <= _GEN_34146;
      end
    end else begin
      rob_uop_28_src1_value <= _GEN_29728;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_28_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1c == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_28_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_28_alu_sel <= _GEN_34466;
        end
      end else begin
        rob_uop_28_alu_sel <= _GEN_34466;
      end
    end else begin
      rob_uop_28_alu_sel <= _GEN_30048;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_29_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1d == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_29_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_29_pc <= _GEN_32739;
        end
      end else begin
        rob_uop_29_pc <= _GEN_32739;
      end
    end else begin
      rob_uop_29_pc <= _GEN_28321;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_29_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1d == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_29_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_29_inst <= _GEN_32803;
        end
      end else begin
        rob_uop_29_inst <= _GEN_32803;
      end
    end else begin
      rob_uop_29_inst <= _GEN_28385;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_29_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1d == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_29_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_29_func_code <= _GEN_32867;
        end
      end else begin
        rob_uop_29_func_code <= _GEN_32867;
      end
    end else begin
      rob_uop_29_func_code <= _GEN_28449;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_29_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1d == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_29_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_29_phy_dst <= _GEN_33251;
        end
      end else begin
        rob_uop_29_phy_dst <= _GEN_33251;
      end
    end else begin
      rob_uop_29_phy_dst <= _GEN_28833;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_29_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1d == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_29_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_29_stale_dst <= _GEN_33315;
        end
      end else begin
        rob_uop_29_stale_dst <= _GEN_33315;
      end
    end else begin
      rob_uop_29_stale_dst <= _GEN_28897;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_29_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1d == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_29_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_29_arch_dst <= _GEN_33379;
        end
      end else begin
        rob_uop_29_arch_dst <= _GEN_33379;
      end
    end else begin
      rob_uop_29_arch_dst <= _GEN_28961;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_29_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1d == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_29_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_29_dst_value <= _GEN_34083;
        end
      end else begin
        rob_uop_29_dst_value <= _GEN_34083;
      end
    end else begin
      rob_uop_29_dst_value <= _GEN_29665;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_29_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1d == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_29_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_29_src1_value <= _GEN_34147;
        end
      end else begin
        rob_uop_29_src1_value <= _GEN_34147;
      end
    end else begin
      rob_uop_29_src1_value <= _GEN_29729;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_29_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1d == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_29_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_29_alu_sel <= _GEN_34467;
        end
      end else begin
        rob_uop_29_alu_sel <= _GEN_34467;
      end
    end else begin
      rob_uop_29_alu_sel <= _GEN_30049;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_30_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1e == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_30_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_30_pc <= _GEN_32740;
        end
      end else begin
        rob_uop_30_pc <= _GEN_32740;
      end
    end else begin
      rob_uop_30_pc <= _GEN_28322;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_30_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1e == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_30_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_30_inst <= _GEN_32804;
        end
      end else begin
        rob_uop_30_inst <= _GEN_32804;
      end
    end else begin
      rob_uop_30_inst <= _GEN_28386;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_30_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1e == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_30_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_30_func_code <= _GEN_32868;
        end
      end else begin
        rob_uop_30_func_code <= _GEN_32868;
      end
    end else begin
      rob_uop_30_func_code <= _GEN_28450;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_30_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1e == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_30_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_30_phy_dst <= _GEN_33252;
        end
      end else begin
        rob_uop_30_phy_dst <= _GEN_33252;
      end
    end else begin
      rob_uop_30_phy_dst <= _GEN_28834;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_30_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1e == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_30_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_30_stale_dst <= _GEN_33316;
        end
      end else begin
        rob_uop_30_stale_dst <= _GEN_33316;
      end
    end else begin
      rob_uop_30_stale_dst <= _GEN_28898;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_30_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1e == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_30_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_30_arch_dst <= _GEN_33380;
        end
      end else begin
        rob_uop_30_arch_dst <= _GEN_33380;
      end
    end else begin
      rob_uop_30_arch_dst <= _GEN_28962;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_30_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1e == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_30_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_30_dst_value <= _GEN_34084;
        end
      end else begin
        rob_uop_30_dst_value <= _GEN_34084;
      end
    end else begin
      rob_uop_30_dst_value <= _GEN_29666;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_30_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1e == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_30_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_30_src1_value <= _GEN_34148;
        end
      end else begin
        rob_uop_30_src1_value <= _GEN_34148;
      end
    end else begin
      rob_uop_30_src1_value <= _GEN_29730;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_30_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1e == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_30_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_30_alu_sel <= _GEN_34468;
        end
      end else begin
        rob_uop_30_alu_sel <= _GEN_34468;
      end
    end else begin
      rob_uop_30_alu_sel <= _GEN_30050;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_31_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1f == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_31_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_31_pc <= _GEN_32741;
        end
      end else begin
        rob_uop_31_pc <= _GEN_32741;
      end
    end else begin
      rob_uop_31_pc <= _GEN_28323;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_31_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1f == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_31_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_31_inst <= _GEN_32805;
        end
      end else begin
        rob_uop_31_inst <= _GEN_32805;
      end
    end else begin
      rob_uop_31_inst <= _GEN_28387;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_31_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1f == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_31_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_31_func_code <= _GEN_32869;
        end
      end else begin
        rob_uop_31_func_code <= _GEN_32869;
      end
    end else begin
      rob_uop_31_func_code <= _GEN_28451;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_31_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1f == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_31_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_31_phy_dst <= _GEN_33253;
        end
      end else begin
        rob_uop_31_phy_dst <= _GEN_33253;
      end
    end else begin
      rob_uop_31_phy_dst <= _GEN_28835;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_31_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1f == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_31_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_31_stale_dst <= _GEN_33317;
        end
      end else begin
        rob_uop_31_stale_dst <= _GEN_33317;
      end
    end else begin
      rob_uop_31_stale_dst <= _GEN_28899;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_31_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1f == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_31_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_31_arch_dst <= _GEN_33381;
        end
      end else begin
        rob_uop_31_arch_dst <= _GEN_33381;
      end
    end else begin
      rob_uop_31_arch_dst <= _GEN_28963;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_31_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1f == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_31_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_31_dst_value <= _GEN_34085;
        end
      end else begin
        rob_uop_31_dst_value <= _GEN_34085;
      end
    end else begin
      rob_uop_31_dst_value <= _GEN_29667;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_31_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1f == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_31_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_31_src1_value <= _GEN_34149;
        end
      end else begin
        rob_uop_31_src1_value <= _GEN_34149;
      end
    end else begin
      rob_uop_31_src1_value <= _GEN_29731;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_31_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h1f == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_31_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_31_alu_sel <= _GEN_34469;
        end
      end else begin
        rob_uop_31_alu_sel <= _GEN_34469;
      end
    end else begin
      rob_uop_31_alu_sel <= _GEN_30051;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_32_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h20 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_32_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_32_pc <= _GEN_32742;
        end
      end else begin
        rob_uop_32_pc <= _GEN_32742;
      end
    end else begin
      rob_uop_32_pc <= _GEN_28324;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_32_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h20 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_32_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_32_inst <= _GEN_32806;
        end
      end else begin
        rob_uop_32_inst <= _GEN_32806;
      end
    end else begin
      rob_uop_32_inst <= _GEN_28388;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_32_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h20 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_32_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_32_func_code <= _GEN_32870;
        end
      end else begin
        rob_uop_32_func_code <= _GEN_32870;
      end
    end else begin
      rob_uop_32_func_code <= _GEN_28452;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_32_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h20 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_32_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_32_phy_dst <= _GEN_33254;
        end
      end else begin
        rob_uop_32_phy_dst <= _GEN_33254;
      end
    end else begin
      rob_uop_32_phy_dst <= _GEN_28836;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_32_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h20 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_32_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_32_stale_dst <= _GEN_33318;
        end
      end else begin
        rob_uop_32_stale_dst <= _GEN_33318;
      end
    end else begin
      rob_uop_32_stale_dst <= _GEN_28900;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_32_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h20 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_32_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_32_arch_dst <= _GEN_33382;
        end
      end else begin
        rob_uop_32_arch_dst <= _GEN_33382;
      end
    end else begin
      rob_uop_32_arch_dst <= _GEN_28964;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_32_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h20 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_32_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_32_dst_value <= _GEN_34086;
        end
      end else begin
        rob_uop_32_dst_value <= _GEN_34086;
      end
    end else begin
      rob_uop_32_dst_value <= _GEN_29668;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_32_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h20 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_32_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_32_src1_value <= _GEN_34150;
        end
      end else begin
        rob_uop_32_src1_value <= _GEN_34150;
      end
    end else begin
      rob_uop_32_src1_value <= _GEN_29732;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_32_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h20 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_32_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_32_alu_sel <= _GEN_34470;
        end
      end else begin
        rob_uop_32_alu_sel <= _GEN_34470;
      end
    end else begin
      rob_uop_32_alu_sel <= _GEN_30052;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_33_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h21 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_33_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_33_pc <= _GEN_32743;
        end
      end else begin
        rob_uop_33_pc <= _GEN_32743;
      end
    end else begin
      rob_uop_33_pc <= _GEN_28325;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_33_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h21 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_33_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_33_inst <= _GEN_32807;
        end
      end else begin
        rob_uop_33_inst <= _GEN_32807;
      end
    end else begin
      rob_uop_33_inst <= _GEN_28389;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_33_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h21 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_33_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_33_func_code <= _GEN_32871;
        end
      end else begin
        rob_uop_33_func_code <= _GEN_32871;
      end
    end else begin
      rob_uop_33_func_code <= _GEN_28453;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_33_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h21 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_33_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_33_phy_dst <= _GEN_33255;
        end
      end else begin
        rob_uop_33_phy_dst <= _GEN_33255;
      end
    end else begin
      rob_uop_33_phy_dst <= _GEN_28837;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_33_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h21 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_33_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_33_stale_dst <= _GEN_33319;
        end
      end else begin
        rob_uop_33_stale_dst <= _GEN_33319;
      end
    end else begin
      rob_uop_33_stale_dst <= _GEN_28901;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_33_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h21 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_33_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_33_arch_dst <= _GEN_33383;
        end
      end else begin
        rob_uop_33_arch_dst <= _GEN_33383;
      end
    end else begin
      rob_uop_33_arch_dst <= _GEN_28965;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_33_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h21 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_33_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_33_dst_value <= _GEN_34087;
        end
      end else begin
        rob_uop_33_dst_value <= _GEN_34087;
      end
    end else begin
      rob_uop_33_dst_value <= _GEN_29669;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_33_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h21 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_33_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_33_src1_value <= _GEN_34151;
        end
      end else begin
        rob_uop_33_src1_value <= _GEN_34151;
      end
    end else begin
      rob_uop_33_src1_value <= _GEN_29733;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_33_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h21 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_33_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_33_alu_sel <= _GEN_34471;
        end
      end else begin
        rob_uop_33_alu_sel <= _GEN_34471;
      end
    end else begin
      rob_uop_33_alu_sel <= _GEN_30053;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_34_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h22 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_34_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_34_pc <= _GEN_32744;
        end
      end else begin
        rob_uop_34_pc <= _GEN_32744;
      end
    end else begin
      rob_uop_34_pc <= _GEN_28326;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_34_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h22 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_34_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_34_inst <= _GEN_32808;
        end
      end else begin
        rob_uop_34_inst <= _GEN_32808;
      end
    end else begin
      rob_uop_34_inst <= _GEN_28390;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_34_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h22 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_34_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_34_func_code <= _GEN_32872;
        end
      end else begin
        rob_uop_34_func_code <= _GEN_32872;
      end
    end else begin
      rob_uop_34_func_code <= _GEN_28454;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_34_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h22 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_34_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_34_phy_dst <= _GEN_33256;
        end
      end else begin
        rob_uop_34_phy_dst <= _GEN_33256;
      end
    end else begin
      rob_uop_34_phy_dst <= _GEN_28838;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_34_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h22 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_34_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_34_stale_dst <= _GEN_33320;
        end
      end else begin
        rob_uop_34_stale_dst <= _GEN_33320;
      end
    end else begin
      rob_uop_34_stale_dst <= _GEN_28902;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_34_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h22 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_34_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_34_arch_dst <= _GEN_33384;
        end
      end else begin
        rob_uop_34_arch_dst <= _GEN_33384;
      end
    end else begin
      rob_uop_34_arch_dst <= _GEN_28966;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_34_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h22 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_34_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_34_dst_value <= _GEN_34088;
        end
      end else begin
        rob_uop_34_dst_value <= _GEN_34088;
      end
    end else begin
      rob_uop_34_dst_value <= _GEN_29670;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_34_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h22 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_34_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_34_src1_value <= _GEN_34152;
        end
      end else begin
        rob_uop_34_src1_value <= _GEN_34152;
      end
    end else begin
      rob_uop_34_src1_value <= _GEN_29734;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_34_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h22 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_34_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_34_alu_sel <= _GEN_34472;
        end
      end else begin
        rob_uop_34_alu_sel <= _GEN_34472;
      end
    end else begin
      rob_uop_34_alu_sel <= _GEN_30054;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_35_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h23 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_35_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_35_pc <= _GEN_32745;
        end
      end else begin
        rob_uop_35_pc <= _GEN_32745;
      end
    end else begin
      rob_uop_35_pc <= _GEN_28327;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_35_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h23 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_35_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_35_inst <= _GEN_32809;
        end
      end else begin
        rob_uop_35_inst <= _GEN_32809;
      end
    end else begin
      rob_uop_35_inst <= _GEN_28391;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_35_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h23 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_35_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_35_func_code <= _GEN_32873;
        end
      end else begin
        rob_uop_35_func_code <= _GEN_32873;
      end
    end else begin
      rob_uop_35_func_code <= _GEN_28455;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_35_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h23 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_35_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_35_phy_dst <= _GEN_33257;
        end
      end else begin
        rob_uop_35_phy_dst <= _GEN_33257;
      end
    end else begin
      rob_uop_35_phy_dst <= _GEN_28839;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_35_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h23 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_35_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_35_stale_dst <= _GEN_33321;
        end
      end else begin
        rob_uop_35_stale_dst <= _GEN_33321;
      end
    end else begin
      rob_uop_35_stale_dst <= _GEN_28903;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_35_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h23 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_35_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_35_arch_dst <= _GEN_33385;
        end
      end else begin
        rob_uop_35_arch_dst <= _GEN_33385;
      end
    end else begin
      rob_uop_35_arch_dst <= _GEN_28967;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_35_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h23 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_35_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_35_dst_value <= _GEN_34089;
        end
      end else begin
        rob_uop_35_dst_value <= _GEN_34089;
      end
    end else begin
      rob_uop_35_dst_value <= _GEN_29671;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_35_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h23 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_35_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_35_src1_value <= _GEN_34153;
        end
      end else begin
        rob_uop_35_src1_value <= _GEN_34153;
      end
    end else begin
      rob_uop_35_src1_value <= _GEN_29735;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_35_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h23 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_35_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_35_alu_sel <= _GEN_34473;
        end
      end else begin
        rob_uop_35_alu_sel <= _GEN_34473;
      end
    end else begin
      rob_uop_35_alu_sel <= _GEN_30055;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_36_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h24 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_36_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_36_pc <= _GEN_32746;
        end
      end else begin
        rob_uop_36_pc <= _GEN_32746;
      end
    end else begin
      rob_uop_36_pc <= _GEN_28328;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_36_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h24 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_36_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_36_inst <= _GEN_32810;
        end
      end else begin
        rob_uop_36_inst <= _GEN_32810;
      end
    end else begin
      rob_uop_36_inst <= _GEN_28392;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_36_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h24 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_36_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_36_func_code <= _GEN_32874;
        end
      end else begin
        rob_uop_36_func_code <= _GEN_32874;
      end
    end else begin
      rob_uop_36_func_code <= _GEN_28456;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_36_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h24 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_36_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_36_phy_dst <= _GEN_33258;
        end
      end else begin
        rob_uop_36_phy_dst <= _GEN_33258;
      end
    end else begin
      rob_uop_36_phy_dst <= _GEN_28840;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_36_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h24 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_36_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_36_stale_dst <= _GEN_33322;
        end
      end else begin
        rob_uop_36_stale_dst <= _GEN_33322;
      end
    end else begin
      rob_uop_36_stale_dst <= _GEN_28904;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_36_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h24 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_36_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_36_arch_dst <= _GEN_33386;
        end
      end else begin
        rob_uop_36_arch_dst <= _GEN_33386;
      end
    end else begin
      rob_uop_36_arch_dst <= _GEN_28968;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_36_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h24 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_36_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_36_dst_value <= _GEN_34090;
        end
      end else begin
        rob_uop_36_dst_value <= _GEN_34090;
      end
    end else begin
      rob_uop_36_dst_value <= _GEN_29672;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_36_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h24 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_36_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_36_src1_value <= _GEN_34154;
        end
      end else begin
        rob_uop_36_src1_value <= _GEN_34154;
      end
    end else begin
      rob_uop_36_src1_value <= _GEN_29736;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_36_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h24 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_36_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_36_alu_sel <= _GEN_34474;
        end
      end else begin
        rob_uop_36_alu_sel <= _GEN_34474;
      end
    end else begin
      rob_uop_36_alu_sel <= _GEN_30056;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_37_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h25 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_37_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_37_pc <= _GEN_32747;
        end
      end else begin
        rob_uop_37_pc <= _GEN_32747;
      end
    end else begin
      rob_uop_37_pc <= _GEN_28329;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_37_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h25 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_37_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_37_inst <= _GEN_32811;
        end
      end else begin
        rob_uop_37_inst <= _GEN_32811;
      end
    end else begin
      rob_uop_37_inst <= _GEN_28393;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_37_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h25 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_37_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_37_func_code <= _GEN_32875;
        end
      end else begin
        rob_uop_37_func_code <= _GEN_32875;
      end
    end else begin
      rob_uop_37_func_code <= _GEN_28457;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_37_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h25 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_37_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_37_phy_dst <= _GEN_33259;
        end
      end else begin
        rob_uop_37_phy_dst <= _GEN_33259;
      end
    end else begin
      rob_uop_37_phy_dst <= _GEN_28841;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_37_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h25 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_37_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_37_stale_dst <= _GEN_33323;
        end
      end else begin
        rob_uop_37_stale_dst <= _GEN_33323;
      end
    end else begin
      rob_uop_37_stale_dst <= _GEN_28905;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_37_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h25 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_37_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_37_arch_dst <= _GEN_33387;
        end
      end else begin
        rob_uop_37_arch_dst <= _GEN_33387;
      end
    end else begin
      rob_uop_37_arch_dst <= _GEN_28969;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_37_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h25 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_37_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_37_dst_value <= _GEN_34091;
        end
      end else begin
        rob_uop_37_dst_value <= _GEN_34091;
      end
    end else begin
      rob_uop_37_dst_value <= _GEN_29673;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_37_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h25 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_37_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_37_src1_value <= _GEN_34155;
        end
      end else begin
        rob_uop_37_src1_value <= _GEN_34155;
      end
    end else begin
      rob_uop_37_src1_value <= _GEN_29737;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_37_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h25 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_37_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_37_alu_sel <= _GEN_34475;
        end
      end else begin
        rob_uop_37_alu_sel <= _GEN_34475;
      end
    end else begin
      rob_uop_37_alu_sel <= _GEN_30057;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_38_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h26 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_38_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_38_pc <= _GEN_32748;
        end
      end else begin
        rob_uop_38_pc <= _GEN_32748;
      end
    end else begin
      rob_uop_38_pc <= _GEN_28330;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_38_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h26 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_38_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_38_inst <= _GEN_32812;
        end
      end else begin
        rob_uop_38_inst <= _GEN_32812;
      end
    end else begin
      rob_uop_38_inst <= _GEN_28394;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_38_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h26 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_38_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_38_func_code <= _GEN_32876;
        end
      end else begin
        rob_uop_38_func_code <= _GEN_32876;
      end
    end else begin
      rob_uop_38_func_code <= _GEN_28458;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_38_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h26 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_38_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_38_phy_dst <= _GEN_33260;
        end
      end else begin
        rob_uop_38_phy_dst <= _GEN_33260;
      end
    end else begin
      rob_uop_38_phy_dst <= _GEN_28842;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_38_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h26 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_38_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_38_stale_dst <= _GEN_33324;
        end
      end else begin
        rob_uop_38_stale_dst <= _GEN_33324;
      end
    end else begin
      rob_uop_38_stale_dst <= _GEN_28906;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_38_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h26 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_38_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_38_arch_dst <= _GEN_33388;
        end
      end else begin
        rob_uop_38_arch_dst <= _GEN_33388;
      end
    end else begin
      rob_uop_38_arch_dst <= _GEN_28970;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_38_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h26 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_38_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_38_dst_value <= _GEN_34092;
        end
      end else begin
        rob_uop_38_dst_value <= _GEN_34092;
      end
    end else begin
      rob_uop_38_dst_value <= _GEN_29674;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_38_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h26 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_38_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_38_src1_value <= _GEN_34156;
        end
      end else begin
        rob_uop_38_src1_value <= _GEN_34156;
      end
    end else begin
      rob_uop_38_src1_value <= _GEN_29738;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_38_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h26 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_38_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_38_alu_sel <= _GEN_34476;
        end
      end else begin
        rob_uop_38_alu_sel <= _GEN_34476;
      end
    end else begin
      rob_uop_38_alu_sel <= _GEN_30058;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_39_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h27 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_39_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_39_pc <= _GEN_32749;
        end
      end else begin
        rob_uop_39_pc <= _GEN_32749;
      end
    end else begin
      rob_uop_39_pc <= _GEN_28331;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_39_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h27 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_39_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_39_inst <= _GEN_32813;
        end
      end else begin
        rob_uop_39_inst <= _GEN_32813;
      end
    end else begin
      rob_uop_39_inst <= _GEN_28395;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_39_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h27 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_39_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_39_func_code <= _GEN_32877;
        end
      end else begin
        rob_uop_39_func_code <= _GEN_32877;
      end
    end else begin
      rob_uop_39_func_code <= _GEN_28459;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_39_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h27 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_39_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_39_phy_dst <= _GEN_33261;
        end
      end else begin
        rob_uop_39_phy_dst <= _GEN_33261;
      end
    end else begin
      rob_uop_39_phy_dst <= _GEN_28843;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_39_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h27 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_39_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_39_stale_dst <= _GEN_33325;
        end
      end else begin
        rob_uop_39_stale_dst <= _GEN_33325;
      end
    end else begin
      rob_uop_39_stale_dst <= _GEN_28907;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_39_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h27 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_39_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_39_arch_dst <= _GEN_33389;
        end
      end else begin
        rob_uop_39_arch_dst <= _GEN_33389;
      end
    end else begin
      rob_uop_39_arch_dst <= _GEN_28971;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_39_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h27 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_39_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_39_dst_value <= _GEN_34093;
        end
      end else begin
        rob_uop_39_dst_value <= _GEN_34093;
      end
    end else begin
      rob_uop_39_dst_value <= _GEN_29675;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_39_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h27 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_39_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_39_src1_value <= _GEN_34157;
        end
      end else begin
        rob_uop_39_src1_value <= _GEN_34157;
      end
    end else begin
      rob_uop_39_src1_value <= _GEN_29739;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_39_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h27 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_39_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_39_alu_sel <= _GEN_34477;
        end
      end else begin
        rob_uop_39_alu_sel <= _GEN_34477;
      end
    end else begin
      rob_uop_39_alu_sel <= _GEN_30059;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_40_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h28 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_40_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_40_pc <= _GEN_32750;
        end
      end else begin
        rob_uop_40_pc <= _GEN_32750;
      end
    end else begin
      rob_uop_40_pc <= _GEN_28332;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_40_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h28 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_40_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_40_inst <= _GEN_32814;
        end
      end else begin
        rob_uop_40_inst <= _GEN_32814;
      end
    end else begin
      rob_uop_40_inst <= _GEN_28396;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_40_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h28 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_40_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_40_func_code <= _GEN_32878;
        end
      end else begin
        rob_uop_40_func_code <= _GEN_32878;
      end
    end else begin
      rob_uop_40_func_code <= _GEN_28460;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_40_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h28 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_40_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_40_phy_dst <= _GEN_33262;
        end
      end else begin
        rob_uop_40_phy_dst <= _GEN_33262;
      end
    end else begin
      rob_uop_40_phy_dst <= _GEN_28844;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_40_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h28 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_40_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_40_stale_dst <= _GEN_33326;
        end
      end else begin
        rob_uop_40_stale_dst <= _GEN_33326;
      end
    end else begin
      rob_uop_40_stale_dst <= _GEN_28908;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_40_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h28 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_40_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_40_arch_dst <= _GEN_33390;
        end
      end else begin
        rob_uop_40_arch_dst <= _GEN_33390;
      end
    end else begin
      rob_uop_40_arch_dst <= _GEN_28972;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_40_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h28 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_40_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_40_dst_value <= _GEN_34094;
        end
      end else begin
        rob_uop_40_dst_value <= _GEN_34094;
      end
    end else begin
      rob_uop_40_dst_value <= _GEN_29676;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_40_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h28 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_40_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_40_src1_value <= _GEN_34158;
        end
      end else begin
        rob_uop_40_src1_value <= _GEN_34158;
      end
    end else begin
      rob_uop_40_src1_value <= _GEN_29740;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_40_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h28 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_40_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_40_alu_sel <= _GEN_34478;
        end
      end else begin
        rob_uop_40_alu_sel <= _GEN_34478;
      end
    end else begin
      rob_uop_40_alu_sel <= _GEN_30060;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_41_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h29 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_41_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_41_pc <= _GEN_32751;
        end
      end else begin
        rob_uop_41_pc <= _GEN_32751;
      end
    end else begin
      rob_uop_41_pc <= _GEN_28333;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_41_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h29 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_41_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_41_inst <= _GEN_32815;
        end
      end else begin
        rob_uop_41_inst <= _GEN_32815;
      end
    end else begin
      rob_uop_41_inst <= _GEN_28397;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_41_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h29 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_41_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_41_func_code <= _GEN_32879;
        end
      end else begin
        rob_uop_41_func_code <= _GEN_32879;
      end
    end else begin
      rob_uop_41_func_code <= _GEN_28461;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_41_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h29 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_41_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_41_phy_dst <= _GEN_33263;
        end
      end else begin
        rob_uop_41_phy_dst <= _GEN_33263;
      end
    end else begin
      rob_uop_41_phy_dst <= _GEN_28845;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_41_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h29 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_41_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_41_stale_dst <= _GEN_33327;
        end
      end else begin
        rob_uop_41_stale_dst <= _GEN_33327;
      end
    end else begin
      rob_uop_41_stale_dst <= _GEN_28909;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_41_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h29 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_41_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_41_arch_dst <= _GEN_33391;
        end
      end else begin
        rob_uop_41_arch_dst <= _GEN_33391;
      end
    end else begin
      rob_uop_41_arch_dst <= _GEN_28973;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_41_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h29 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_41_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_41_dst_value <= _GEN_34095;
        end
      end else begin
        rob_uop_41_dst_value <= _GEN_34095;
      end
    end else begin
      rob_uop_41_dst_value <= _GEN_29677;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_41_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h29 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_41_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_41_src1_value <= _GEN_34159;
        end
      end else begin
        rob_uop_41_src1_value <= _GEN_34159;
      end
    end else begin
      rob_uop_41_src1_value <= _GEN_29741;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_41_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h29 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_41_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_41_alu_sel <= _GEN_34479;
        end
      end else begin
        rob_uop_41_alu_sel <= _GEN_34479;
      end
    end else begin
      rob_uop_41_alu_sel <= _GEN_30061;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_42_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2a == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_42_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_42_pc <= _GEN_32752;
        end
      end else begin
        rob_uop_42_pc <= _GEN_32752;
      end
    end else begin
      rob_uop_42_pc <= _GEN_28334;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_42_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2a == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_42_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_42_inst <= _GEN_32816;
        end
      end else begin
        rob_uop_42_inst <= _GEN_32816;
      end
    end else begin
      rob_uop_42_inst <= _GEN_28398;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_42_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2a == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_42_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_42_func_code <= _GEN_32880;
        end
      end else begin
        rob_uop_42_func_code <= _GEN_32880;
      end
    end else begin
      rob_uop_42_func_code <= _GEN_28462;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_42_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2a == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_42_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_42_phy_dst <= _GEN_33264;
        end
      end else begin
        rob_uop_42_phy_dst <= _GEN_33264;
      end
    end else begin
      rob_uop_42_phy_dst <= _GEN_28846;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_42_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2a == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_42_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_42_stale_dst <= _GEN_33328;
        end
      end else begin
        rob_uop_42_stale_dst <= _GEN_33328;
      end
    end else begin
      rob_uop_42_stale_dst <= _GEN_28910;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_42_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2a == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_42_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_42_arch_dst <= _GEN_33392;
        end
      end else begin
        rob_uop_42_arch_dst <= _GEN_33392;
      end
    end else begin
      rob_uop_42_arch_dst <= _GEN_28974;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_42_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2a == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_42_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_42_dst_value <= _GEN_34096;
        end
      end else begin
        rob_uop_42_dst_value <= _GEN_34096;
      end
    end else begin
      rob_uop_42_dst_value <= _GEN_29678;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_42_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2a == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_42_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_42_src1_value <= _GEN_34160;
        end
      end else begin
        rob_uop_42_src1_value <= _GEN_34160;
      end
    end else begin
      rob_uop_42_src1_value <= _GEN_29742;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_42_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2a == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_42_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_42_alu_sel <= _GEN_34480;
        end
      end else begin
        rob_uop_42_alu_sel <= _GEN_34480;
      end
    end else begin
      rob_uop_42_alu_sel <= _GEN_30062;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_43_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2b == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_43_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_43_pc <= _GEN_32753;
        end
      end else begin
        rob_uop_43_pc <= _GEN_32753;
      end
    end else begin
      rob_uop_43_pc <= _GEN_28335;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_43_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2b == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_43_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_43_inst <= _GEN_32817;
        end
      end else begin
        rob_uop_43_inst <= _GEN_32817;
      end
    end else begin
      rob_uop_43_inst <= _GEN_28399;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_43_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2b == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_43_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_43_func_code <= _GEN_32881;
        end
      end else begin
        rob_uop_43_func_code <= _GEN_32881;
      end
    end else begin
      rob_uop_43_func_code <= _GEN_28463;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_43_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2b == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_43_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_43_phy_dst <= _GEN_33265;
        end
      end else begin
        rob_uop_43_phy_dst <= _GEN_33265;
      end
    end else begin
      rob_uop_43_phy_dst <= _GEN_28847;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_43_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2b == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_43_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_43_stale_dst <= _GEN_33329;
        end
      end else begin
        rob_uop_43_stale_dst <= _GEN_33329;
      end
    end else begin
      rob_uop_43_stale_dst <= _GEN_28911;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_43_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2b == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_43_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_43_arch_dst <= _GEN_33393;
        end
      end else begin
        rob_uop_43_arch_dst <= _GEN_33393;
      end
    end else begin
      rob_uop_43_arch_dst <= _GEN_28975;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_43_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2b == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_43_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_43_dst_value <= _GEN_34097;
        end
      end else begin
        rob_uop_43_dst_value <= _GEN_34097;
      end
    end else begin
      rob_uop_43_dst_value <= _GEN_29679;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_43_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2b == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_43_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_43_src1_value <= _GEN_34161;
        end
      end else begin
        rob_uop_43_src1_value <= _GEN_34161;
      end
    end else begin
      rob_uop_43_src1_value <= _GEN_29743;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_43_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2b == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_43_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_43_alu_sel <= _GEN_34481;
        end
      end else begin
        rob_uop_43_alu_sel <= _GEN_34481;
      end
    end else begin
      rob_uop_43_alu_sel <= _GEN_30063;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_44_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2c == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_44_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_44_pc <= _GEN_32754;
        end
      end else begin
        rob_uop_44_pc <= _GEN_32754;
      end
    end else begin
      rob_uop_44_pc <= _GEN_28336;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_44_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2c == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_44_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_44_inst <= _GEN_32818;
        end
      end else begin
        rob_uop_44_inst <= _GEN_32818;
      end
    end else begin
      rob_uop_44_inst <= _GEN_28400;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_44_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2c == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_44_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_44_func_code <= _GEN_32882;
        end
      end else begin
        rob_uop_44_func_code <= _GEN_32882;
      end
    end else begin
      rob_uop_44_func_code <= _GEN_28464;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_44_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2c == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_44_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_44_phy_dst <= _GEN_33266;
        end
      end else begin
        rob_uop_44_phy_dst <= _GEN_33266;
      end
    end else begin
      rob_uop_44_phy_dst <= _GEN_28848;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_44_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2c == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_44_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_44_stale_dst <= _GEN_33330;
        end
      end else begin
        rob_uop_44_stale_dst <= _GEN_33330;
      end
    end else begin
      rob_uop_44_stale_dst <= _GEN_28912;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_44_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2c == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_44_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_44_arch_dst <= _GEN_33394;
        end
      end else begin
        rob_uop_44_arch_dst <= _GEN_33394;
      end
    end else begin
      rob_uop_44_arch_dst <= _GEN_28976;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_44_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2c == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_44_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_44_dst_value <= _GEN_34098;
        end
      end else begin
        rob_uop_44_dst_value <= _GEN_34098;
      end
    end else begin
      rob_uop_44_dst_value <= _GEN_29680;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_44_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2c == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_44_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_44_src1_value <= _GEN_34162;
        end
      end else begin
        rob_uop_44_src1_value <= _GEN_34162;
      end
    end else begin
      rob_uop_44_src1_value <= _GEN_29744;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_44_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2c == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_44_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_44_alu_sel <= _GEN_34482;
        end
      end else begin
        rob_uop_44_alu_sel <= _GEN_34482;
      end
    end else begin
      rob_uop_44_alu_sel <= _GEN_30064;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_45_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2d == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_45_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_45_pc <= _GEN_32755;
        end
      end else begin
        rob_uop_45_pc <= _GEN_32755;
      end
    end else begin
      rob_uop_45_pc <= _GEN_28337;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_45_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2d == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_45_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_45_inst <= _GEN_32819;
        end
      end else begin
        rob_uop_45_inst <= _GEN_32819;
      end
    end else begin
      rob_uop_45_inst <= _GEN_28401;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_45_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2d == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_45_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_45_func_code <= _GEN_32883;
        end
      end else begin
        rob_uop_45_func_code <= _GEN_32883;
      end
    end else begin
      rob_uop_45_func_code <= _GEN_28465;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_45_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2d == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_45_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_45_phy_dst <= _GEN_33267;
        end
      end else begin
        rob_uop_45_phy_dst <= _GEN_33267;
      end
    end else begin
      rob_uop_45_phy_dst <= _GEN_28849;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_45_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2d == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_45_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_45_stale_dst <= _GEN_33331;
        end
      end else begin
        rob_uop_45_stale_dst <= _GEN_33331;
      end
    end else begin
      rob_uop_45_stale_dst <= _GEN_28913;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_45_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2d == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_45_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_45_arch_dst <= _GEN_33395;
        end
      end else begin
        rob_uop_45_arch_dst <= _GEN_33395;
      end
    end else begin
      rob_uop_45_arch_dst <= _GEN_28977;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_45_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2d == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_45_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_45_dst_value <= _GEN_34099;
        end
      end else begin
        rob_uop_45_dst_value <= _GEN_34099;
      end
    end else begin
      rob_uop_45_dst_value <= _GEN_29681;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_45_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2d == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_45_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_45_src1_value <= _GEN_34163;
        end
      end else begin
        rob_uop_45_src1_value <= _GEN_34163;
      end
    end else begin
      rob_uop_45_src1_value <= _GEN_29745;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_45_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2d == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_45_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_45_alu_sel <= _GEN_34483;
        end
      end else begin
        rob_uop_45_alu_sel <= _GEN_34483;
      end
    end else begin
      rob_uop_45_alu_sel <= _GEN_30065;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_46_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2e == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_46_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_46_pc <= _GEN_32756;
        end
      end else begin
        rob_uop_46_pc <= _GEN_32756;
      end
    end else begin
      rob_uop_46_pc <= _GEN_28338;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_46_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2e == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_46_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_46_inst <= _GEN_32820;
        end
      end else begin
        rob_uop_46_inst <= _GEN_32820;
      end
    end else begin
      rob_uop_46_inst <= _GEN_28402;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_46_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2e == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_46_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_46_func_code <= _GEN_32884;
        end
      end else begin
        rob_uop_46_func_code <= _GEN_32884;
      end
    end else begin
      rob_uop_46_func_code <= _GEN_28466;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_46_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2e == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_46_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_46_phy_dst <= _GEN_33268;
        end
      end else begin
        rob_uop_46_phy_dst <= _GEN_33268;
      end
    end else begin
      rob_uop_46_phy_dst <= _GEN_28850;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_46_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2e == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_46_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_46_stale_dst <= _GEN_33332;
        end
      end else begin
        rob_uop_46_stale_dst <= _GEN_33332;
      end
    end else begin
      rob_uop_46_stale_dst <= _GEN_28914;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_46_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2e == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_46_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_46_arch_dst <= _GEN_33396;
        end
      end else begin
        rob_uop_46_arch_dst <= _GEN_33396;
      end
    end else begin
      rob_uop_46_arch_dst <= _GEN_28978;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_46_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2e == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_46_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_46_dst_value <= _GEN_34100;
        end
      end else begin
        rob_uop_46_dst_value <= _GEN_34100;
      end
    end else begin
      rob_uop_46_dst_value <= _GEN_29682;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_46_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2e == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_46_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_46_src1_value <= _GEN_34164;
        end
      end else begin
        rob_uop_46_src1_value <= _GEN_34164;
      end
    end else begin
      rob_uop_46_src1_value <= _GEN_29746;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_46_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2e == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_46_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_46_alu_sel <= _GEN_34484;
        end
      end else begin
        rob_uop_46_alu_sel <= _GEN_34484;
      end
    end else begin
      rob_uop_46_alu_sel <= _GEN_30066;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_47_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2f == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_47_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_47_pc <= _GEN_32757;
        end
      end else begin
        rob_uop_47_pc <= _GEN_32757;
      end
    end else begin
      rob_uop_47_pc <= _GEN_28339;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_47_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2f == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_47_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_47_inst <= _GEN_32821;
        end
      end else begin
        rob_uop_47_inst <= _GEN_32821;
      end
    end else begin
      rob_uop_47_inst <= _GEN_28403;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_47_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2f == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_47_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_47_func_code <= _GEN_32885;
        end
      end else begin
        rob_uop_47_func_code <= _GEN_32885;
      end
    end else begin
      rob_uop_47_func_code <= _GEN_28467;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_47_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2f == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_47_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_47_phy_dst <= _GEN_33269;
        end
      end else begin
        rob_uop_47_phy_dst <= _GEN_33269;
      end
    end else begin
      rob_uop_47_phy_dst <= _GEN_28851;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_47_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2f == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_47_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_47_stale_dst <= _GEN_33333;
        end
      end else begin
        rob_uop_47_stale_dst <= _GEN_33333;
      end
    end else begin
      rob_uop_47_stale_dst <= _GEN_28915;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_47_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2f == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_47_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_47_arch_dst <= _GEN_33397;
        end
      end else begin
        rob_uop_47_arch_dst <= _GEN_33397;
      end
    end else begin
      rob_uop_47_arch_dst <= _GEN_28979;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_47_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2f == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_47_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_47_dst_value <= _GEN_34101;
        end
      end else begin
        rob_uop_47_dst_value <= _GEN_34101;
      end
    end else begin
      rob_uop_47_dst_value <= _GEN_29683;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_47_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2f == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_47_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_47_src1_value <= _GEN_34165;
        end
      end else begin
        rob_uop_47_src1_value <= _GEN_34165;
      end
    end else begin
      rob_uop_47_src1_value <= _GEN_29747;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_47_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h2f == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_47_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_47_alu_sel <= _GEN_34485;
        end
      end else begin
        rob_uop_47_alu_sel <= _GEN_34485;
      end
    end else begin
      rob_uop_47_alu_sel <= _GEN_30067;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_48_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h30 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_48_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_48_pc <= _GEN_32758;
        end
      end else begin
        rob_uop_48_pc <= _GEN_32758;
      end
    end else begin
      rob_uop_48_pc <= _GEN_28340;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_48_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h30 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_48_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_48_inst <= _GEN_32822;
        end
      end else begin
        rob_uop_48_inst <= _GEN_32822;
      end
    end else begin
      rob_uop_48_inst <= _GEN_28404;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_48_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h30 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_48_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_48_func_code <= _GEN_32886;
        end
      end else begin
        rob_uop_48_func_code <= _GEN_32886;
      end
    end else begin
      rob_uop_48_func_code <= _GEN_28468;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_48_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h30 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_48_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_48_phy_dst <= _GEN_33270;
        end
      end else begin
        rob_uop_48_phy_dst <= _GEN_33270;
      end
    end else begin
      rob_uop_48_phy_dst <= _GEN_28852;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_48_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h30 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_48_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_48_stale_dst <= _GEN_33334;
        end
      end else begin
        rob_uop_48_stale_dst <= _GEN_33334;
      end
    end else begin
      rob_uop_48_stale_dst <= _GEN_28916;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_48_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h30 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_48_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_48_arch_dst <= _GEN_33398;
        end
      end else begin
        rob_uop_48_arch_dst <= _GEN_33398;
      end
    end else begin
      rob_uop_48_arch_dst <= _GEN_28980;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_48_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h30 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_48_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_48_dst_value <= _GEN_34102;
        end
      end else begin
        rob_uop_48_dst_value <= _GEN_34102;
      end
    end else begin
      rob_uop_48_dst_value <= _GEN_29684;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_48_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h30 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_48_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_48_src1_value <= _GEN_34166;
        end
      end else begin
        rob_uop_48_src1_value <= _GEN_34166;
      end
    end else begin
      rob_uop_48_src1_value <= _GEN_29748;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_48_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h30 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_48_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_48_alu_sel <= _GEN_34486;
        end
      end else begin
        rob_uop_48_alu_sel <= _GEN_34486;
      end
    end else begin
      rob_uop_48_alu_sel <= _GEN_30068;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_49_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h31 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_49_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_49_pc <= _GEN_32759;
        end
      end else begin
        rob_uop_49_pc <= _GEN_32759;
      end
    end else begin
      rob_uop_49_pc <= _GEN_28341;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_49_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h31 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_49_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_49_inst <= _GEN_32823;
        end
      end else begin
        rob_uop_49_inst <= _GEN_32823;
      end
    end else begin
      rob_uop_49_inst <= _GEN_28405;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_49_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h31 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_49_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_49_func_code <= _GEN_32887;
        end
      end else begin
        rob_uop_49_func_code <= _GEN_32887;
      end
    end else begin
      rob_uop_49_func_code <= _GEN_28469;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_49_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h31 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_49_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_49_phy_dst <= _GEN_33271;
        end
      end else begin
        rob_uop_49_phy_dst <= _GEN_33271;
      end
    end else begin
      rob_uop_49_phy_dst <= _GEN_28853;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_49_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h31 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_49_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_49_stale_dst <= _GEN_33335;
        end
      end else begin
        rob_uop_49_stale_dst <= _GEN_33335;
      end
    end else begin
      rob_uop_49_stale_dst <= _GEN_28917;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_49_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h31 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_49_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_49_arch_dst <= _GEN_33399;
        end
      end else begin
        rob_uop_49_arch_dst <= _GEN_33399;
      end
    end else begin
      rob_uop_49_arch_dst <= _GEN_28981;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_49_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h31 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_49_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_49_dst_value <= _GEN_34103;
        end
      end else begin
        rob_uop_49_dst_value <= _GEN_34103;
      end
    end else begin
      rob_uop_49_dst_value <= _GEN_29685;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_49_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h31 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_49_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_49_src1_value <= _GEN_34167;
        end
      end else begin
        rob_uop_49_src1_value <= _GEN_34167;
      end
    end else begin
      rob_uop_49_src1_value <= _GEN_29749;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_49_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h31 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_49_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_49_alu_sel <= _GEN_34487;
        end
      end else begin
        rob_uop_49_alu_sel <= _GEN_34487;
      end
    end else begin
      rob_uop_49_alu_sel <= _GEN_30069;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_50_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h32 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_50_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_50_pc <= _GEN_32760;
        end
      end else begin
        rob_uop_50_pc <= _GEN_32760;
      end
    end else begin
      rob_uop_50_pc <= _GEN_28342;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_50_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h32 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_50_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_50_inst <= _GEN_32824;
        end
      end else begin
        rob_uop_50_inst <= _GEN_32824;
      end
    end else begin
      rob_uop_50_inst <= _GEN_28406;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_50_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h32 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_50_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_50_func_code <= _GEN_32888;
        end
      end else begin
        rob_uop_50_func_code <= _GEN_32888;
      end
    end else begin
      rob_uop_50_func_code <= _GEN_28470;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_50_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h32 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_50_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_50_phy_dst <= _GEN_33272;
        end
      end else begin
        rob_uop_50_phy_dst <= _GEN_33272;
      end
    end else begin
      rob_uop_50_phy_dst <= _GEN_28854;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_50_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h32 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_50_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_50_stale_dst <= _GEN_33336;
        end
      end else begin
        rob_uop_50_stale_dst <= _GEN_33336;
      end
    end else begin
      rob_uop_50_stale_dst <= _GEN_28918;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_50_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h32 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_50_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_50_arch_dst <= _GEN_33400;
        end
      end else begin
        rob_uop_50_arch_dst <= _GEN_33400;
      end
    end else begin
      rob_uop_50_arch_dst <= _GEN_28982;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_50_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h32 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_50_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_50_dst_value <= _GEN_34104;
        end
      end else begin
        rob_uop_50_dst_value <= _GEN_34104;
      end
    end else begin
      rob_uop_50_dst_value <= _GEN_29686;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_50_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h32 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_50_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_50_src1_value <= _GEN_34168;
        end
      end else begin
        rob_uop_50_src1_value <= _GEN_34168;
      end
    end else begin
      rob_uop_50_src1_value <= _GEN_29750;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_50_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h32 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_50_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_50_alu_sel <= _GEN_34488;
        end
      end else begin
        rob_uop_50_alu_sel <= _GEN_34488;
      end
    end else begin
      rob_uop_50_alu_sel <= _GEN_30070;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_51_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h33 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_51_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_51_pc <= _GEN_32761;
        end
      end else begin
        rob_uop_51_pc <= _GEN_32761;
      end
    end else begin
      rob_uop_51_pc <= _GEN_28343;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_51_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h33 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_51_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_51_inst <= _GEN_32825;
        end
      end else begin
        rob_uop_51_inst <= _GEN_32825;
      end
    end else begin
      rob_uop_51_inst <= _GEN_28407;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_51_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h33 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_51_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_51_func_code <= _GEN_32889;
        end
      end else begin
        rob_uop_51_func_code <= _GEN_32889;
      end
    end else begin
      rob_uop_51_func_code <= _GEN_28471;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_51_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h33 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_51_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_51_phy_dst <= _GEN_33273;
        end
      end else begin
        rob_uop_51_phy_dst <= _GEN_33273;
      end
    end else begin
      rob_uop_51_phy_dst <= _GEN_28855;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_51_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h33 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_51_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_51_stale_dst <= _GEN_33337;
        end
      end else begin
        rob_uop_51_stale_dst <= _GEN_33337;
      end
    end else begin
      rob_uop_51_stale_dst <= _GEN_28919;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_51_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h33 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_51_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_51_arch_dst <= _GEN_33401;
        end
      end else begin
        rob_uop_51_arch_dst <= _GEN_33401;
      end
    end else begin
      rob_uop_51_arch_dst <= _GEN_28983;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_51_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h33 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_51_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_51_dst_value <= _GEN_34105;
        end
      end else begin
        rob_uop_51_dst_value <= _GEN_34105;
      end
    end else begin
      rob_uop_51_dst_value <= _GEN_29687;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_51_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h33 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_51_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_51_src1_value <= _GEN_34169;
        end
      end else begin
        rob_uop_51_src1_value <= _GEN_34169;
      end
    end else begin
      rob_uop_51_src1_value <= _GEN_29751;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_51_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h33 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_51_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_51_alu_sel <= _GEN_34489;
        end
      end else begin
        rob_uop_51_alu_sel <= _GEN_34489;
      end
    end else begin
      rob_uop_51_alu_sel <= _GEN_30071;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_52_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h34 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_52_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_52_pc <= _GEN_32762;
        end
      end else begin
        rob_uop_52_pc <= _GEN_32762;
      end
    end else begin
      rob_uop_52_pc <= _GEN_28344;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_52_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h34 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_52_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_52_inst <= _GEN_32826;
        end
      end else begin
        rob_uop_52_inst <= _GEN_32826;
      end
    end else begin
      rob_uop_52_inst <= _GEN_28408;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_52_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h34 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_52_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_52_func_code <= _GEN_32890;
        end
      end else begin
        rob_uop_52_func_code <= _GEN_32890;
      end
    end else begin
      rob_uop_52_func_code <= _GEN_28472;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_52_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h34 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_52_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_52_phy_dst <= _GEN_33274;
        end
      end else begin
        rob_uop_52_phy_dst <= _GEN_33274;
      end
    end else begin
      rob_uop_52_phy_dst <= _GEN_28856;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_52_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h34 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_52_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_52_stale_dst <= _GEN_33338;
        end
      end else begin
        rob_uop_52_stale_dst <= _GEN_33338;
      end
    end else begin
      rob_uop_52_stale_dst <= _GEN_28920;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_52_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h34 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_52_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_52_arch_dst <= _GEN_33402;
        end
      end else begin
        rob_uop_52_arch_dst <= _GEN_33402;
      end
    end else begin
      rob_uop_52_arch_dst <= _GEN_28984;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_52_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h34 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_52_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_52_dst_value <= _GEN_34106;
        end
      end else begin
        rob_uop_52_dst_value <= _GEN_34106;
      end
    end else begin
      rob_uop_52_dst_value <= _GEN_29688;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_52_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h34 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_52_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_52_src1_value <= _GEN_34170;
        end
      end else begin
        rob_uop_52_src1_value <= _GEN_34170;
      end
    end else begin
      rob_uop_52_src1_value <= _GEN_29752;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_52_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h34 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_52_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_52_alu_sel <= _GEN_34490;
        end
      end else begin
        rob_uop_52_alu_sel <= _GEN_34490;
      end
    end else begin
      rob_uop_52_alu_sel <= _GEN_30072;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_53_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h35 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_53_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_53_pc <= _GEN_32763;
        end
      end else begin
        rob_uop_53_pc <= _GEN_32763;
      end
    end else begin
      rob_uop_53_pc <= _GEN_28345;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_53_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h35 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_53_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_53_inst <= _GEN_32827;
        end
      end else begin
        rob_uop_53_inst <= _GEN_32827;
      end
    end else begin
      rob_uop_53_inst <= _GEN_28409;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_53_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h35 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_53_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_53_func_code <= _GEN_32891;
        end
      end else begin
        rob_uop_53_func_code <= _GEN_32891;
      end
    end else begin
      rob_uop_53_func_code <= _GEN_28473;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_53_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h35 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_53_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_53_phy_dst <= _GEN_33275;
        end
      end else begin
        rob_uop_53_phy_dst <= _GEN_33275;
      end
    end else begin
      rob_uop_53_phy_dst <= _GEN_28857;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_53_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h35 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_53_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_53_stale_dst <= _GEN_33339;
        end
      end else begin
        rob_uop_53_stale_dst <= _GEN_33339;
      end
    end else begin
      rob_uop_53_stale_dst <= _GEN_28921;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_53_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h35 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_53_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_53_arch_dst <= _GEN_33403;
        end
      end else begin
        rob_uop_53_arch_dst <= _GEN_33403;
      end
    end else begin
      rob_uop_53_arch_dst <= _GEN_28985;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_53_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h35 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_53_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_53_dst_value <= _GEN_34107;
        end
      end else begin
        rob_uop_53_dst_value <= _GEN_34107;
      end
    end else begin
      rob_uop_53_dst_value <= _GEN_29689;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_53_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h35 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_53_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_53_src1_value <= _GEN_34171;
        end
      end else begin
        rob_uop_53_src1_value <= _GEN_34171;
      end
    end else begin
      rob_uop_53_src1_value <= _GEN_29753;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_53_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h35 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_53_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_53_alu_sel <= _GEN_34491;
        end
      end else begin
        rob_uop_53_alu_sel <= _GEN_34491;
      end
    end else begin
      rob_uop_53_alu_sel <= _GEN_30073;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_54_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h36 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_54_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_54_pc <= _GEN_32764;
        end
      end else begin
        rob_uop_54_pc <= _GEN_32764;
      end
    end else begin
      rob_uop_54_pc <= _GEN_28346;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_54_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h36 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_54_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_54_inst <= _GEN_32828;
        end
      end else begin
        rob_uop_54_inst <= _GEN_32828;
      end
    end else begin
      rob_uop_54_inst <= _GEN_28410;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_54_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h36 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_54_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_54_func_code <= _GEN_32892;
        end
      end else begin
        rob_uop_54_func_code <= _GEN_32892;
      end
    end else begin
      rob_uop_54_func_code <= _GEN_28474;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_54_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h36 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_54_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_54_phy_dst <= _GEN_33276;
        end
      end else begin
        rob_uop_54_phy_dst <= _GEN_33276;
      end
    end else begin
      rob_uop_54_phy_dst <= _GEN_28858;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_54_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h36 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_54_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_54_stale_dst <= _GEN_33340;
        end
      end else begin
        rob_uop_54_stale_dst <= _GEN_33340;
      end
    end else begin
      rob_uop_54_stale_dst <= _GEN_28922;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_54_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h36 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_54_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_54_arch_dst <= _GEN_33404;
        end
      end else begin
        rob_uop_54_arch_dst <= _GEN_33404;
      end
    end else begin
      rob_uop_54_arch_dst <= _GEN_28986;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_54_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h36 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_54_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_54_dst_value <= _GEN_34108;
        end
      end else begin
        rob_uop_54_dst_value <= _GEN_34108;
      end
    end else begin
      rob_uop_54_dst_value <= _GEN_29690;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_54_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h36 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_54_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_54_src1_value <= _GEN_34172;
        end
      end else begin
        rob_uop_54_src1_value <= _GEN_34172;
      end
    end else begin
      rob_uop_54_src1_value <= _GEN_29754;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_54_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h36 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_54_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_54_alu_sel <= _GEN_34492;
        end
      end else begin
        rob_uop_54_alu_sel <= _GEN_34492;
      end
    end else begin
      rob_uop_54_alu_sel <= _GEN_30074;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_55_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h37 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_55_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_55_pc <= _GEN_32765;
        end
      end else begin
        rob_uop_55_pc <= _GEN_32765;
      end
    end else begin
      rob_uop_55_pc <= _GEN_28347;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_55_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h37 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_55_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_55_inst <= _GEN_32829;
        end
      end else begin
        rob_uop_55_inst <= _GEN_32829;
      end
    end else begin
      rob_uop_55_inst <= _GEN_28411;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_55_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h37 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_55_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_55_func_code <= _GEN_32893;
        end
      end else begin
        rob_uop_55_func_code <= _GEN_32893;
      end
    end else begin
      rob_uop_55_func_code <= _GEN_28475;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_55_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h37 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_55_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_55_phy_dst <= _GEN_33277;
        end
      end else begin
        rob_uop_55_phy_dst <= _GEN_33277;
      end
    end else begin
      rob_uop_55_phy_dst <= _GEN_28859;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_55_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h37 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_55_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_55_stale_dst <= _GEN_33341;
        end
      end else begin
        rob_uop_55_stale_dst <= _GEN_33341;
      end
    end else begin
      rob_uop_55_stale_dst <= _GEN_28923;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_55_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h37 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_55_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_55_arch_dst <= _GEN_33405;
        end
      end else begin
        rob_uop_55_arch_dst <= _GEN_33405;
      end
    end else begin
      rob_uop_55_arch_dst <= _GEN_28987;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_55_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h37 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_55_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_55_dst_value <= _GEN_34109;
        end
      end else begin
        rob_uop_55_dst_value <= _GEN_34109;
      end
    end else begin
      rob_uop_55_dst_value <= _GEN_29691;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_55_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h37 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_55_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_55_src1_value <= _GEN_34173;
        end
      end else begin
        rob_uop_55_src1_value <= _GEN_34173;
      end
    end else begin
      rob_uop_55_src1_value <= _GEN_29755;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_55_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h37 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_55_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_55_alu_sel <= _GEN_34493;
        end
      end else begin
        rob_uop_55_alu_sel <= _GEN_34493;
      end
    end else begin
      rob_uop_55_alu_sel <= _GEN_30075;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_56_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h38 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_56_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_56_pc <= _GEN_32766;
        end
      end else begin
        rob_uop_56_pc <= _GEN_32766;
      end
    end else begin
      rob_uop_56_pc <= _GEN_28348;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_56_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h38 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_56_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_56_inst <= _GEN_32830;
        end
      end else begin
        rob_uop_56_inst <= _GEN_32830;
      end
    end else begin
      rob_uop_56_inst <= _GEN_28412;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_56_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h38 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_56_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_56_func_code <= _GEN_32894;
        end
      end else begin
        rob_uop_56_func_code <= _GEN_32894;
      end
    end else begin
      rob_uop_56_func_code <= _GEN_28476;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_56_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h38 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_56_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_56_phy_dst <= _GEN_33278;
        end
      end else begin
        rob_uop_56_phy_dst <= _GEN_33278;
      end
    end else begin
      rob_uop_56_phy_dst <= _GEN_28860;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_56_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h38 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_56_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_56_stale_dst <= _GEN_33342;
        end
      end else begin
        rob_uop_56_stale_dst <= _GEN_33342;
      end
    end else begin
      rob_uop_56_stale_dst <= _GEN_28924;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_56_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h38 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_56_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_56_arch_dst <= _GEN_33406;
        end
      end else begin
        rob_uop_56_arch_dst <= _GEN_33406;
      end
    end else begin
      rob_uop_56_arch_dst <= _GEN_28988;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_56_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h38 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_56_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_56_dst_value <= _GEN_34110;
        end
      end else begin
        rob_uop_56_dst_value <= _GEN_34110;
      end
    end else begin
      rob_uop_56_dst_value <= _GEN_29692;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_56_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h38 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_56_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_56_src1_value <= _GEN_34174;
        end
      end else begin
        rob_uop_56_src1_value <= _GEN_34174;
      end
    end else begin
      rob_uop_56_src1_value <= _GEN_29756;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_56_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h38 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_56_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_56_alu_sel <= _GEN_34494;
        end
      end else begin
        rob_uop_56_alu_sel <= _GEN_34494;
      end
    end else begin
      rob_uop_56_alu_sel <= _GEN_30076;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_57_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h39 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_57_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_57_pc <= _GEN_32767;
        end
      end else begin
        rob_uop_57_pc <= _GEN_32767;
      end
    end else begin
      rob_uop_57_pc <= _GEN_28349;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_57_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h39 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_57_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_57_inst <= _GEN_32831;
        end
      end else begin
        rob_uop_57_inst <= _GEN_32831;
      end
    end else begin
      rob_uop_57_inst <= _GEN_28413;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_57_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h39 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_57_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_57_func_code <= _GEN_32895;
        end
      end else begin
        rob_uop_57_func_code <= _GEN_32895;
      end
    end else begin
      rob_uop_57_func_code <= _GEN_28477;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_57_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h39 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_57_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_57_phy_dst <= _GEN_33279;
        end
      end else begin
        rob_uop_57_phy_dst <= _GEN_33279;
      end
    end else begin
      rob_uop_57_phy_dst <= _GEN_28861;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_57_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h39 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_57_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_57_stale_dst <= _GEN_33343;
        end
      end else begin
        rob_uop_57_stale_dst <= _GEN_33343;
      end
    end else begin
      rob_uop_57_stale_dst <= _GEN_28925;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_57_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h39 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_57_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_57_arch_dst <= _GEN_33407;
        end
      end else begin
        rob_uop_57_arch_dst <= _GEN_33407;
      end
    end else begin
      rob_uop_57_arch_dst <= _GEN_28989;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_57_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h39 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_57_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_57_dst_value <= _GEN_34111;
        end
      end else begin
        rob_uop_57_dst_value <= _GEN_34111;
      end
    end else begin
      rob_uop_57_dst_value <= _GEN_29693;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_57_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h39 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_57_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_57_src1_value <= _GEN_34175;
        end
      end else begin
        rob_uop_57_src1_value <= _GEN_34175;
      end
    end else begin
      rob_uop_57_src1_value <= _GEN_29757;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_57_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h39 == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_57_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_57_alu_sel <= _GEN_34495;
        end
      end else begin
        rob_uop_57_alu_sel <= _GEN_34495;
      end
    end else begin
      rob_uop_57_alu_sel <= _GEN_30077;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_58_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3a == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_58_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_58_pc <= _GEN_32768;
        end
      end else begin
        rob_uop_58_pc <= _GEN_32768;
      end
    end else begin
      rob_uop_58_pc <= _GEN_28350;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_58_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3a == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_58_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_58_inst <= _GEN_32832;
        end
      end else begin
        rob_uop_58_inst <= _GEN_32832;
      end
    end else begin
      rob_uop_58_inst <= _GEN_28414;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_58_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3a == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_58_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_58_func_code <= _GEN_32896;
        end
      end else begin
        rob_uop_58_func_code <= _GEN_32896;
      end
    end else begin
      rob_uop_58_func_code <= _GEN_28478;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_58_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3a == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_58_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_58_phy_dst <= _GEN_33280;
        end
      end else begin
        rob_uop_58_phy_dst <= _GEN_33280;
      end
    end else begin
      rob_uop_58_phy_dst <= _GEN_28862;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_58_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3a == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_58_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_58_stale_dst <= _GEN_33344;
        end
      end else begin
        rob_uop_58_stale_dst <= _GEN_33344;
      end
    end else begin
      rob_uop_58_stale_dst <= _GEN_28926;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_58_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3a == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_58_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_58_arch_dst <= _GEN_33408;
        end
      end else begin
        rob_uop_58_arch_dst <= _GEN_33408;
      end
    end else begin
      rob_uop_58_arch_dst <= _GEN_28990;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_58_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3a == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_58_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_58_dst_value <= _GEN_34112;
        end
      end else begin
        rob_uop_58_dst_value <= _GEN_34112;
      end
    end else begin
      rob_uop_58_dst_value <= _GEN_29694;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_58_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3a == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_58_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_58_src1_value <= _GEN_34176;
        end
      end else begin
        rob_uop_58_src1_value <= _GEN_34176;
      end
    end else begin
      rob_uop_58_src1_value <= _GEN_29758;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_58_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3a == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_58_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_58_alu_sel <= _GEN_34496;
        end
      end else begin
        rob_uop_58_alu_sel <= _GEN_34496;
      end
    end else begin
      rob_uop_58_alu_sel <= _GEN_30078;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_59_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3b == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_59_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_59_pc <= _GEN_32769;
        end
      end else begin
        rob_uop_59_pc <= _GEN_32769;
      end
    end else begin
      rob_uop_59_pc <= _GEN_28351;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_59_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3b == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_59_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_59_inst <= _GEN_32833;
        end
      end else begin
        rob_uop_59_inst <= _GEN_32833;
      end
    end else begin
      rob_uop_59_inst <= _GEN_28415;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_59_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3b == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_59_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_59_func_code <= _GEN_32897;
        end
      end else begin
        rob_uop_59_func_code <= _GEN_32897;
      end
    end else begin
      rob_uop_59_func_code <= _GEN_28479;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_59_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3b == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_59_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_59_phy_dst <= _GEN_33281;
        end
      end else begin
        rob_uop_59_phy_dst <= _GEN_33281;
      end
    end else begin
      rob_uop_59_phy_dst <= _GEN_28863;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_59_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3b == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_59_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_59_stale_dst <= _GEN_33345;
        end
      end else begin
        rob_uop_59_stale_dst <= _GEN_33345;
      end
    end else begin
      rob_uop_59_stale_dst <= _GEN_28927;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_59_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3b == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_59_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_59_arch_dst <= _GEN_33409;
        end
      end else begin
        rob_uop_59_arch_dst <= _GEN_33409;
      end
    end else begin
      rob_uop_59_arch_dst <= _GEN_28991;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_59_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3b == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_59_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_59_dst_value <= _GEN_34113;
        end
      end else begin
        rob_uop_59_dst_value <= _GEN_34113;
      end
    end else begin
      rob_uop_59_dst_value <= _GEN_29695;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_59_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3b == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_59_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_59_src1_value <= _GEN_34177;
        end
      end else begin
        rob_uop_59_src1_value <= _GEN_34177;
      end
    end else begin
      rob_uop_59_src1_value <= _GEN_29759;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_59_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3b == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_59_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_59_alu_sel <= _GEN_34497;
        end
      end else begin
        rob_uop_59_alu_sel <= _GEN_34497;
      end
    end else begin
      rob_uop_59_alu_sel <= _GEN_30079;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_60_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3c == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_60_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_60_pc <= _GEN_32770;
        end
      end else begin
        rob_uop_60_pc <= _GEN_32770;
      end
    end else begin
      rob_uop_60_pc <= _GEN_28352;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_60_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3c == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_60_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_60_inst <= _GEN_32834;
        end
      end else begin
        rob_uop_60_inst <= _GEN_32834;
      end
    end else begin
      rob_uop_60_inst <= _GEN_28416;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_60_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3c == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_60_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_60_func_code <= _GEN_32898;
        end
      end else begin
        rob_uop_60_func_code <= _GEN_32898;
      end
    end else begin
      rob_uop_60_func_code <= _GEN_28480;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_60_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3c == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_60_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_60_phy_dst <= _GEN_33282;
        end
      end else begin
        rob_uop_60_phy_dst <= _GEN_33282;
      end
    end else begin
      rob_uop_60_phy_dst <= _GEN_28864;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_60_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3c == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_60_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_60_stale_dst <= _GEN_33346;
        end
      end else begin
        rob_uop_60_stale_dst <= _GEN_33346;
      end
    end else begin
      rob_uop_60_stale_dst <= _GEN_28928;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_60_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3c == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_60_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_60_arch_dst <= _GEN_33410;
        end
      end else begin
        rob_uop_60_arch_dst <= _GEN_33410;
      end
    end else begin
      rob_uop_60_arch_dst <= _GEN_28992;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_60_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3c == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_60_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_60_dst_value <= _GEN_34114;
        end
      end else begin
        rob_uop_60_dst_value <= _GEN_34114;
      end
    end else begin
      rob_uop_60_dst_value <= _GEN_29696;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_60_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3c == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_60_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_60_src1_value <= _GEN_34178;
        end
      end else begin
        rob_uop_60_src1_value <= _GEN_34178;
      end
    end else begin
      rob_uop_60_src1_value <= _GEN_29760;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_60_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3c == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_60_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_60_alu_sel <= _GEN_34498;
        end
      end else begin
        rob_uop_60_alu_sel <= _GEN_34498;
      end
    end else begin
      rob_uop_60_alu_sel <= _GEN_30080;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_61_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3d == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_61_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_61_pc <= _GEN_32771;
        end
      end else begin
        rob_uop_61_pc <= _GEN_32771;
      end
    end else begin
      rob_uop_61_pc <= _GEN_28353;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_61_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3d == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_61_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_61_inst <= _GEN_32835;
        end
      end else begin
        rob_uop_61_inst <= _GEN_32835;
      end
    end else begin
      rob_uop_61_inst <= _GEN_28417;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_61_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3d == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_61_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_61_func_code <= _GEN_32899;
        end
      end else begin
        rob_uop_61_func_code <= _GEN_32899;
      end
    end else begin
      rob_uop_61_func_code <= _GEN_28481;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_61_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3d == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_61_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_61_phy_dst <= _GEN_33283;
        end
      end else begin
        rob_uop_61_phy_dst <= _GEN_33283;
      end
    end else begin
      rob_uop_61_phy_dst <= _GEN_28865;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_61_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3d == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_61_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_61_stale_dst <= _GEN_33347;
        end
      end else begin
        rob_uop_61_stale_dst <= _GEN_33347;
      end
    end else begin
      rob_uop_61_stale_dst <= _GEN_28929;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_61_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3d == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_61_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_61_arch_dst <= _GEN_33411;
        end
      end else begin
        rob_uop_61_arch_dst <= _GEN_33411;
      end
    end else begin
      rob_uop_61_arch_dst <= _GEN_28993;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_61_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3d == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_61_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_61_dst_value <= _GEN_34115;
        end
      end else begin
        rob_uop_61_dst_value <= _GEN_34115;
      end
    end else begin
      rob_uop_61_dst_value <= _GEN_29697;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_61_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3d == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_61_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_61_src1_value <= _GEN_34179;
        end
      end else begin
        rob_uop_61_src1_value <= _GEN_34179;
      end
    end else begin
      rob_uop_61_src1_value <= _GEN_29761;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_61_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3d == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_61_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_61_alu_sel <= _GEN_34499;
        end
      end else begin
        rob_uop_61_alu_sel <= _GEN_34499;
      end
    end else begin
      rob_uop_61_alu_sel <= _GEN_30081;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_62_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3e == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_62_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_62_pc <= _GEN_32772;
        end
      end else begin
        rob_uop_62_pc <= _GEN_32772;
      end
    end else begin
      rob_uop_62_pc <= _GEN_28354;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_62_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3e == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_62_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_62_inst <= _GEN_32836;
        end
      end else begin
        rob_uop_62_inst <= _GEN_32836;
      end
    end else begin
      rob_uop_62_inst <= _GEN_28418;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_62_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3e == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_62_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_62_func_code <= _GEN_32900;
        end
      end else begin
        rob_uop_62_func_code <= _GEN_32900;
      end
    end else begin
      rob_uop_62_func_code <= _GEN_28482;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_62_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3e == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_62_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_62_phy_dst <= _GEN_33284;
        end
      end else begin
        rob_uop_62_phy_dst <= _GEN_33284;
      end
    end else begin
      rob_uop_62_phy_dst <= _GEN_28866;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_62_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3e == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_62_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_62_stale_dst <= _GEN_33348;
        end
      end else begin
        rob_uop_62_stale_dst <= _GEN_33348;
      end
    end else begin
      rob_uop_62_stale_dst <= _GEN_28930;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_62_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3e == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_62_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_62_arch_dst <= _GEN_33412;
        end
      end else begin
        rob_uop_62_arch_dst <= _GEN_33412;
      end
    end else begin
      rob_uop_62_arch_dst <= _GEN_28994;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_62_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3e == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_62_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_62_dst_value <= _GEN_34116;
        end
      end else begin
        rob_uop_62_dst_value <= _GEN_34116;
      end
    end else begin
      rob_uop_62_dst_value <= _GEN_29698;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_62_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3e == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_62_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_62_src1_value <= _GEN_34180;
        end
      end else begin
        rob_uop_62_src1_value <= _GEN_34180;
      end
    end else begin
      rob_uop_62_src1_value <= _GEN_29762;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_62_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3e == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_62_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_62_alu_sel <= _GEN_34500;
        end
      end else begin
        rob_uop_62_alu_sel <= _GEN_34500;
      end
    end else begin
      rob_uop_62_alu_sel <= _GEN_30082;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_63_pc <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3f == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_63_pc <= io_i_ex_res_packs_1_uop_pc; // @[rob.scala 174:51]
        end else begin
          rob_uop_63_pc <= _GEN_32773;
        end
      end else begin
        rob_uop_63_pc <= _GEN_32773;
      end
    end else begin
      rob_uop_63_pc <= _GEN_28355;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_63_inst <= 32'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3f == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_63_inst <= io_i_ex_res_packs_1_uop_inst; // @[rob.scala 174:51]
        end else begin
          rob_uop_63_inst <= _GEN_32837;
        end
      end else begin
        rob_uop_63_inst <= _GEN_32837;
      end
    end else begin
      rob_uop_63_inst <= _GEN_28419;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_63_func_code <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3f == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_63_func_code <= io_i_ex_res_packs_1_uop_func_code; // @[rob.scala 174:51]
        end else begin
          rob_uop_63_func_code <= _GEN_32901;
        end
      end else begin
        rob_uop_63_func_code <= _GEN_32901;
      end
    end else begin
      rob_uop_63_func_code <= _GEN_28483;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_63_phy_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3f == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_63_phy_dst <= io_i_ex_res_packs_1_uop_phy_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_63_phy_dst <= _GEN_33285;
        end
      end else begin
        rob_uop_63_phy_dst <= _GEN_33285;
      end
    end else begin
      rob_uop_63_phy_dst <= _GEN_28867;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_63_stale_dst <= 7'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3f == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_63_stale_dst <= io_i_ex_res_packs_1_uop_stale_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_63_stale_dst <= _GEN_33349;
        end
      end else begin
        rob_uop_63_stale_dst <= _GEN_33349;
      end
    end else begin
      rob_uop_63_stale_dst <= _GEN_28931;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_63_arch_dst <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3f == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_63_arch_dst <= io_i_ex_res_packs_1_uop_arch_dst; // @[rob.scala 174:51]
        end else begin
          rob_uop_63_arch_dst <= _GEN_33413;
        end
      end else begin
        rob_uop_63_arch_dst <= _GEN_33413;
      end
    end else begin
      rob_uop_63_arch_dst <= _GEN_28995;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_63_dst_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3f == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_63_dst_value <= io_i_ex_res_packs_1_uop_dst_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_63_dst_value <= _GEN_34117;
        end
      end else begin
        rob_uop_63_dst_value <= _GEN_34117;
      end
    end else begin
      rob_uop_63_dst_value <= _GEN_29699;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_63_src1_value <= 64'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3f == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_63_src1_value <= io_i_ex_res_packs_1_uop_src1_value; // @[rob.scala 174:51]
        end else begin
          rob_uop_63_src1_value <= _GEN_34181;
        end
      end else begin
        rob_uop_63_src1_value <= _GEN_34181;
      end
    end else begin
      rob_uop_63_src1_value <= _GEN_29763;
    end
    if (reset) begin // @[rob.scala 82:26]
      rob_uop_63_alu_sel <= 5'h0; // @[rob.scala 82:26]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        if (6'h3f == io_i_ex_res_packs_1_uop_rob_idx[5:0]) begin // @[rob.scala 174:51]
          rob_uop_63_alu_sel <= io_i_ex_res_packs_1_uop_alu_sel; // @[rob.scala 174:51]
        end else begin
          rob_uop_63_alu_sel <= _GEN_34501;
        end
      end else begin
        rob_uop_63_alu_sel <= _GEN_34501;
      end
    end else begin
      rob_uop_63_alu_sel <= _GEN_30083;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_0 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_0 <= _GEN_36870;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_0 <= _GEN_32518;
      end else begin
        rob_done_0 <= _GEN_30276;
      end
    end else begin
      rob_done_0 <= _GEN_30276;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_1 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_1 <= _GEN_36871;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_1 <= _GEN_32519;
      end else begin
        rob_done_1 <= _GEN_30277;
      end
    end else begin
      rob_done_1 <= _GEN_30277;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_2 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_2 <= _GEN_36872;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_2 <= _GEN_32520;
      end else begin
        rob_done_2 <= _GEN_30278;
      end
    end else begin
      rob_done_2 <= _GEN_30278;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_3 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_3 <= _GEN_36873;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_3 <= _GEN_32521;
      end else begin
        rob_done_3 <= _GEN_30279;
      end
    end else begin
      rob_done_3 <= _GEN_30279;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_4 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_4 <= _GEN_36874;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_4 <= _GEN_32522;
      end else begin
        rob_done_4 <= _GEN_30280;
      end
    end else begin
      rob_done_4 <= _GEN_30280;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_5 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_5 <= _GEN_36875;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_5 <= _GEN_32523;
      end else begin
        rob_done_5 <= _GEN_30281;
      end
    end else begin
      rob_done_5 <= _GEN_30281;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_6 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_6 <= _GEN_36876;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_6 <= _GEN_32524;
      end else begin
        rob_done_6 <= _GEN_30282;
      end
    end else begin
      rob_done_6 <= _GEN_30282;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_7 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_7 <= _GEN_36877;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_7 <= _GEN_32525;
      end else begin
        rob_done_7 <= _GEN_30283;
      end
    end else begin
      rob_done_7 <= _GEN_30283;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_8 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_8 <= _GEN_36878;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_8 <= _GEN_32526;
      end else begin
        rob_done_8 <= _GEN_30284;
      end
    end else begin
      rob_done_8 <= _GEN_30284;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_9 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_9 <= _GEN_36879;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_9 <= _GEN_32527;
      end else begin
        rob_done_9 <= _GEN_30285;
      end
    end else begin
      rob_done_9 <= _GEN_30285;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_10 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_10 <= _GEN_36880;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_10 <= _GEN_32528;
      end else begin
        rob_done_10 <= _GEN_30286;
      end
    end else begin
      rob_done_10 <= _GEN_30286;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_11 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_11 <= _GEN_36881;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_11 <= _GEN_32529;
      end else begin
        rob_done_11 <= _GEN_30287;
      end
    end else begin
      rob_done_11 <= _GEN_30287;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_12 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_12 <= _GEN_36882;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_12 <= _GEN_32530;
      end else begin
        rob_done_12 <= _GEN_30288;
      end
    end else begin
      rob_done_12 <= _GEN_30288;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_13 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_13 <= _GEN_36883;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_13 <= _GEN_32531;
      end else begin
        rob_done_13 <= _GEN_30289;
      end
    end else begin
      rob_done_13 <= _GEN_30289;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_14 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_14 <= _GEN_36884;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_14 <= _GEN_32532;
      end else begin
        rob_done_14 <= _GEN_30290;
      end
    end else begin
      rob_done_14 <= _GEN_30290;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_15 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_15 <= _GEN_36885;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_15 <= _GEN_32533;
      end else begin
        rob_done_15 <= _GEN_30291;
      end
    end else begin
      rob_done_15 <= _GEN_30291;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_16 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_16 <= _GEN_36886;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_16 <= _GEN_32534;
      end else begin
        rob_done_16 <= _GEN_30292;
      end
    end else begin
      rob_done_16 <= _GEN_30292;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_17 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_17 <= _GEN_36887;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_17 <= _GEN_32535;
      end else begin
        rob_done_17 <= _GEN_30293;
      end
    end else begin
      rob_done_17 <= _GEN_30293;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_18 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_18 <= _GEN_36888;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_18 <= _GEN_32536;
      end else begin
        rob_done_18 <= _GEN_30294;
      end
    end else begin
      rob_done_18 <= _GEN_30294;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_19 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_19 <= _GEN_36889;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_19 <= _GEN_32537;
      end else begin
        rob_done_19 <= _GEN_30295;
      end
    end else begin
      rob_done_19 <= _GEN_30295;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_20 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_20 <= _GEN_36890;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_20 <= _GEN_32538;
      end else begin
        rob_done_20 <= _GEN_30296;
      end
    end else begin
      rob_done_20 <= _GEN_30296;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_21 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_21 <= _GEN_36891;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_21 <= _GEN_32539;
      end else begin
        rob_done_21 <= _GEN_30297;
      end
    end else begin
      rob_done_21 <= _GEN_30297;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_22 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_22 <= _GEN_36892;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_22 <= _GEN_32540;
      end else begin
        rob_done_22 <= _GEN_30298;
      end
    end else begin
      rob_done_22 <= _GEN_30298;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_23 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_23 <= _GEN_36893;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_23 <= _GEN_32541;
      end else begin
        rob_done_23 <= _GEN_30299;
      end
    end else begin
      rob_done_23 <= _GEN_30299;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_24 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_24 <= _GEN_36894;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_24 <= _GEN_32542;
      end else begin
        rob_done_24 <= _GEN_30300;
      end
    end else begin
      rob_done_24 <= _GEN_30300;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_25 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_25 <= _GEN_36895;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_25 <= _GEN_32543;
      end else begin
        rob_done_25 <= _GEN_30301;
      end
    end else begin
      rob_done_25 <= _GEN_30301;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_26 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_26 <= _GEN_36896;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_26 <= _GEN_32544;
      end else begin
        rob_done_26 <= _GEN_30302;
      end
    end else begin
      rob_done_26 <= _GEN_30302;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_27 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_27 <= _GEN_36897;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_27 <= _GEN_32545;
      end else begin
        rob_done_27 <= _GEN_30303;
      end
    end else begin
      rob_done_27 <= _GEN_30303;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_28 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_28 <= _GEN_36898;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_28 <= _GEN_32546;
      end else begin
        rob_done_28 <= _GEN_30304;
      end
    end else begin
      rob_done_28 <= _GEN_30304;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_29 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_29 <= _GEN_36899;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_29 <= _GEN_32547;
      end else begin
        rob_done_29 <= _GEN_30305;
      end
    end else begin
      rob_done_29 <= _GEN_30305;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_30 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_30 <= _GEN_36900;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_30 <= _GEN_32548;
      end else begin
        rob_done_30 <= _GEN_30306;
      end
    end else begin
      rob_done_30 <= _GEN_30306;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_31 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_31 <= _GEN_36901;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_31 <= _GEN_32549;
      end else begin
        rob_done_31 <= _GEN_30307;
      end
    end else begin
      rob_done_31 <= _GEN_30307;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_32 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_32 <= _GEN_36902;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_32 <= _GEN_32550;
      end else begin
        rob_done_32 <= _GEN_30308;
      end
    end else begin
      rob_done_32 <= _GEN_30308;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_33 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_33 <= _GEN_36903;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_33 <= _GEN_32551;
      end else begin
        rob_done_33 <= _GEN_30309;
      end
    end else begin
      rob_done_33 <= _GEN_30309;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_34 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_34 <= _GEN_36904;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_34 <= _GEN_32552;
      end else begin
        rob_done_34 <= _GEN_30310;
      end
    end else begin
      rob_done_34 <= _GEN_30310;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_35 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_35 <= _GEN_36905;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_35 <= _GEN_32553;
      end else begin
        rob_done_35 <= _GEN_30311;
      end
    end else begin
      rob_done_35 <= _GEN_30311;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_36 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_36 <= _GEN_36906;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_36 <= _GEN_32554;
      end else begin
        rob_done_36 <= _GEN_30312;
      end
    end else begin
      rob_done_36 <= _GEN_30312;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_37 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_37 <= _GEN_36907;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_37 <= _GEN_32555;
      end else begin
        rob_done_37 <= _GEN_30313;
      end
    end else begin
      rob_done_37 <= _GEN_30313;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_38 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_38 <= _GEN_36908;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_38 <= _GEN_32556;
      end else begin
        rob_done_38 <= _GEN_30314;
      end
    end else begin
      rob_done_38 <= _GEN_30314;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_39 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_39 <= _GEN_36909;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_39 <= _GEN_32557;
      end else begin
        rob_done_39 <= _GEN_30315;
      end
    end else begin
      rob_done_39 <= _GEN_30315;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_40 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_40 <= _GEN_36910;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_40 <= _GEN_32558;
      end else begin
        rob_done_40 <= _GEN_30316;
      end
    end else begin
      rob_done_40 <= _GEN_30316;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_41 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_41 <= _GEN_36911;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_41 <= _GEN_32559;
      end else begin
        rob_done_41 <= _GEN_30317;
      end
    end else begin
      rob_done_41 <= _GEN_30317;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_42 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_42 <= _GEN_36912;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_42 <= _GEN_32560;
      end else begin
        rob_done_42 <= _GEN_30318;
      end
    end else begin
      rob_done_42 <= _GEN_30318;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_43 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_43 <= _GEN_36913;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_43 <= _GEN_32561;
      end else begin
        rob_done_43 <= _GEN_30319;
      end
    end else begin
      rob_done_43 <= _GEN_30319;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_44 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_44 <= _GEN_36914;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_44 <= _GEN_32562;
      end else begin
        rob_done_44 <= _GEN_30320;
      end
    end else begin
      rob_done_44 <= _GEN_30320;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_45 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_45 <= _GEN_36915;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_45 <= _GEN_32563;
      end else begin
        rob_done_45 <= _GEN_30321;
      end
    end else begin
      rob_done_45 <= _GEN_30321;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_46 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_46 <= _GEN_36916;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_46 <= _GEN_32564;
      end else begin
        rob_done_46 <= _GEN_30322;
      end
    end else begin
      rob_done_46 <= _GEN_30322;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_47 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_47 <= _GEN_36917;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_47 <= _GEN_32565;
      end else begin
        rob_done_47 <= _GEN_30323;
      end
    end else begin
      rob_done_47 <= _GEN_30323;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_48 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_48 <= _GEN_36918;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_48 <= _GEN_32566;
      end else begin
        rob_done_48 <= _GEN_30324;
      end
    end else begin
      rob_done_48 <= _GEN_30324;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_49 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_49 <= _GEN_36919;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_49 <= _GEN_32567;
      end else begin
        rob_done_49 <= _GEN_30325;
      end
    end else begin
      rob_done_49 <= _GEN_30325;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_50 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_50 <= _GEN_36920;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_50 <= _GEN_32568;
      end else begin
        rob_done_50 <= _GEN_30326;
      end
    end else begin
      rob_done_50 <= _GEN_30326;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_51 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_51 <= _GEN_36921;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_51 <= _GEN_32569;
      end else begin
        rob_done_51 <= _GEN_30327;
      end
    end else begin
      rob_done_51 <= _GEN_30327;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_52 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_52 <= _GEN_36922;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_52 <= _GEN_32570;
      end else begin
        rob_done_52 <= _GEN_30328;
      end
    end else begin
      rob_done_52 <= _GEN_30328;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_53 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_53 <= _GEN_36923;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_53 <= _GEN_32571;
      end else begin
        rob_done_53 <= _GEN_30329;
      end
    end else begin
      rob_done_53 <= _GEN_30329;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_54 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_54 <= _GEN_36924;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_54 <= _GEN_32572;
      end else begin
        rob_done_54 <= _GEN_30330;
      end
    end else begin
      rob_done_54 <= _GEN_30330;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_55 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_55 <= _GEN_36925;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_55 <= _GEN_32573;
      end else begin
        rob_done_55 <= _GEN_30331;
      end
    end else begin
      rob_done_55 <= _GEN_30331;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_56 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_56 <= _GEN_36926;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_56 <= _GEN_32574;
      end else begin
        rob_done_56 <= _GEN_30332;
      end
    end else begin
      rob_done_56 <= _GEN_30332;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_57 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_57 <= _GEN_36927;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_57 <= _GEN_32575;
      end else begin
        rob_done_57 <= _GEN_30333;
      end
    end else begin
      rob_done_57 <= _GEN_30333;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_58 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_58 <= _GEN_36928;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_58 <= _GEN_32576;
      end else begin
        rob_done_58 <= _GEN_30334;
      end
    end else begin
      rob_done_58 <= _GEN_30334;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_59 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_59 <= _GEN_36929;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_59 <= _GEN_32577;
      end else begin
        rob_done_59 <= _GEN_30335;
      end
    end else begin
      rob_done_59 <= _GEN_30335;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_60 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_60 <= _GEN_36930;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_60 <= _GEN_32578;
      end else begin
        rob_done_60 <= _GEN_30336;
      end
    end else begin
      rob_done_60 <= _GEN_30336;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_61 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_61 <= _GEN_36931;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_61 <= _GEN_32579;
      end else begin
        rob_done_61 <= _GEN_30337;
      end
    end else begin
      rob_done_61 <= _GEN_30337;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_62 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_62 <= _GEN_36932;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_62 <= _GEN_32580;
      end else begin
        rob_done_62 <= _GEN_30338;
      end
    end else begin
      rob_done_62 <= _GEN_30338;
    end
    if (reset) begin // @[rob.scala 84:27]
      rob_done_63 <= 1'h0; // @[rob.scala 84:27]
    end else if (_next_will_commit_0_T_6) begin // @[rob.scala 164:36]
      if (io_i_ex_res_packs_1_valid) begin // @[rob.scala 172:39]
        rob_done_63 <= _GEN_36933;
      end else if (io_i_ex_res_packs_0_valid) begin // @[rob.scala 166:39]
        rob_done_63 <= _GEN_32581;
      end else begin
        rob_done_63 <= _GEN_30339;
      end
    end else begin
      rob_done_63 <= _GEN_30339;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  commit_ptr = _RAND_0[6:0];
  _RAND_1 = {1{`RANDOM}};
  allocate_ptr = _RAND_1[6:0];
  _RAND_2 = {1{`RANDOM}};
  rob_state = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  last_pc_redirect = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  will_commit_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  rob_valid_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  rob_valid_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  rob_valid_2 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  rob_valid_3 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  rob_valid_4 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  rob_valid_5 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  rob_valid_6 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  rob_valid_7 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  rob_valid_8 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  rob_valid_9 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  rob_valid_10 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  rob_valid_11 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  rob_valid_12 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  rob_valid_13 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  rob_valid_14 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  rob_valid_15 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  rob_valid_16 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  rob_valid_17 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  rob_valid_18 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  rob_valid_19 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  rob_valid_20 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  rob_valid_21 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  rob_valid_22 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  rob_valid_23 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  rob_valid_24 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  rob_valid_25 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  rob_valid_26 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  rob_valid_27 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  rob_valid_28 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  rob_valid_29 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  rob_valid_30 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  rob_valid_31 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  rob_valid_32 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  rob_valid_33 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  rob_valid_34 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  rob_valid_35 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  rob_valid_36 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  rob_valid_37 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  rob_valid_38 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  rob_valid_39 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  rob_valid_40 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  rob_valid_41 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  rob_valid_42 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  rob_valid_43 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  rob_valid_44 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  rob_valid_45 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  rob_valid_46 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  rob_valid_47 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  rob_valid_48 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  rob_valid_49 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  rob_valid_50 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  rob_valid_51 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  rob_valid_52 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  rob_valid_53 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  rob_valid_54 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  rob_valid_55 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  rob_valid_56 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  rob_valid_57 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  rob_valid_58 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  rob_valid_59 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  rob_valid_60 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  rob_valid_61 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  rob_valid_62 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  rob_valid_63 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  rob_uop_0_pc = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  rob_uop_0_inst = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  rob_uop_0_func_code = _RAND_71[6:0];
  _RAND_72 = {1{`RANDOM}};
  rob_uop_0_phy_dst = _RAND_72[6:0];
  _RAND_73 = {1{`RANDOM}};
  rob_uop_0_stale_dst = _RAND_73[6:0];
  _RAND_74 = {1{`RANDOM}};
  rob_uop_0_arch_dst = _RAND_74[4:0];
  _RAND_75 = {2{`RANDOM}};
  rob_uop_0_dst_value = _RAND_75[63:0];
  _RAND_76 = {2{`RANDOM}};
  rob_uop_0_src1_value = _RAND_76[63:0];
  _RAND_77 = {1{`RANDOM}};
  rob_uop_0_alu_sel = _RAND_77[4:0];
  _RAND_78 = {1{`RANDOM}};
  rob_uop_1_pc = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  rob_uop_1_inst = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  rob_uop_1_func_code = _RAND_80[6:0];
  _RAND_81 = {1{`RANDOM}};
  rob_uop_1_phy_dst = _RAND_81[6:0];
  _RAND_82 = {1{`RANDOM}};
  rob_uop_1_stale_dst = _RAND_82[6:0];
  _RAND_83 = {1{`RANDOM}};
  rob_uop_1_arch_dst = _RAND_83[4:0];
  _RAND_84 = {2{`RANDOM}};
  rob_uop_1_dst_value = _RAND_84[63:0];
  _RAND_85 = {2{`RANDOM}};
  rob_uop_1_src1_value = _RAND_85[63:0];
  _RAND_86 = {1{`RANDOM}};
  rob_uop_1_alu_sel = _RAND_86[4:0];
  _RAND_87 = {1{`RANDOM}};
  rob_uop_2_pc = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  rob_uop_2_inst = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  rob_uop_2_func_code = _RAND_89[6:0];
  _RAND_90 = {1{`RANDOM}};
  rob_uop_2_phy_dst = _RAND_90[6:0];
  _RAND_91 = {1{`RANDOM}};
  rob_uop_2_stale_dst = _RAND_91[6:0];
  _RAND_92 = {1{`RANDOM}};
  rob_uop_2_arch_dst = _RAND_92[4:0];
  _RAND_93 = {2{`RANDOM}};
  rob_uop_2_dst_value = _RAND_93[63:0];
  _RAND_94 = {2{`RANDOM}};
  rob_uop_2_src1_value = _RAND_94[63:0];
  _RAND_95 = {1{`RANDOM}};
  rob_uop_2_alu_sel = _RAND_95[4:0];
  _RAND_96 = {1{`RANDOM}};
  rob_uop_3_pc = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  rob_uop_3_inst = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  rob_uop_3_func_code = _RAND_98[6:0];
  _RAND_99 = {1{`RANDOM}};
  rob_uop_3_phy_dst = _RAND_99[6:0];
  _RAND_100 = {1{`RANDOM}};
  rob_uop_3_stale_dst = _RAND_100[6:0];
  _RAND_101 = {1{`RANDOM}};
  rob_uop_3_arch_dst = _RAND_101[4:0];
  _RAND_102 = {2{`RANDOM}};
  rob_uop_3_dst_value = _RAND_102[63:0];
  _RAND_103 = {2{`RANDOM}};
  rob_uop_3_src1_value = _RAND_103[63:0];
  _RAND_104 = {1{`RANDOM}};
  rob_uop_3_alu_sel = _RAND_104[4:0];
  _RAND_105 = {1{`RANDOM}};
  rob_uop_4_pc = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  rob_uop_4_inst = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  rob_uop_4_func_code = _RAND_107[6:0];
  _RAND_108 = {1{`RANDOM}};
  rob_uop_4_phy_dst = _RAND_108[6:0];
  _RAND_109 = {1{`RANDOM}};
  rob_uop_4_stale_dst = _RAND_109[6:0];
  _RAND_110 = {1{`RANDOM}};
  rob_uop_4_arch_dst = _RAND_110[4:0];
  _RAND_111 = {2{`RANDOM}};
  rob_uop_4_dst_value = _RAND_111[63:0];
  _RAND_112 = {2{`RANDOM}};
  rob_uop_4_src1_value = _RAND_112[63:0];
  _RAND_113 = {1{`RANDOM}};
  rob_uop_4_alu_sel = _RAND_113[4:0];
  _RAND_114 = {1{`RANDOM}};
  rob_uop_5_pc = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  rob_uop_5_inst = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  rob_uop_5_func_code = _RAND_116[6:0];
  _RAND_117 = {1{`RANDOM}};
  rob_uop_5_phy_dst = _RAND_117[6:0];
  _RAND_118 = {1{`RANDOM}};
  rob_uop_5_stale_dst = _RAND_118[6:0];
  _RAND_119 = {1{`RANDOM}};
  rob_uop_5_arch_dst = _RAND_119[4:0];
  _RAND_120 = {2{`RANDOM}};
  rob_uop_5_dst_value = _RAND_120[63:0];
  _RAND_121 = {2{`RANDOM}};
  rob_uop_5_src1_value = _RAND_121[63:0];
  _RAND_122 = {1{`RANDOM}};
  rob_uop_5_alu_sel = _RAND_122[4:0];
  _RAND_123 = {1{`RANDOM}};
  rob_uop_6_pc = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  rob_uop_6_inst = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  rob_uop_6_func_code = _RAND_125[6:0];
  _RAND_126 = {1{`RANDOM}};
  rob_uop_6_phy_dst = _RAND_126[6:0];
  _RAND_127 = {1{`RANDOM}};
  rob_uop_6_stale_dst = _RAND_127[6:0];
  _RAND_128 = {1{`RANDOM}};
  rob_uop_6_arch_dst = _RAND_128[4:0];
  _RAND_129 = {2{`RANDOM}};
  rob_uop_6_dst_value = _RAND_129[63:0];
  _RAND_130 = {2{`RANDOM}};
  rob_uop_6_src1_value = _RAND_130[63:0];
  _RAND_131 = {1{`RANDOM}};
  rob_uop_6_alu_sel = _RAND_131[4:0];
  _RAND_132 = {1{`RANDOM}};
  rob_uop_7_pc = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  rob_uop_7_inst = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  rob_uop_7_func_code = _RAND_134[6:0];
  _RAND_135 = {1{`RANDOM}};
  rob_uop_7_phy_dst = _RAND_135[6:0];
  _RAND_136 = {1{`RANDOM}};
  rob_uop_7_stale_dst = _RAND_136[6:0];
  _RAND_137 = {1{`RANDOM}};
  rob_uop_7_arch_dst = _RAND_137[4:0];
  _RAND_138 = {2{`RANDOM}};
  rob_uop_7_dst_value = _RAND_138[63:0];
  _RAND_139 = {2{`RANDOM}};
  rob_uop_7_src1_value = _RAND_139[63:0];
  _RAND_140 = {1{`RANDOM}};
  rob_uop_7_alu_sel = _RAND_140[4:0];
  _RAND_141 = {1{`RANDOM}};
  rob_uop_8_pc = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  rob_uop_8_inst = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  rob_uop_8_func_code = _RAND_143[6:0];
  _RAND_144 = {1{`RANDOM}};
  rob_uop_8_phy_dst = _RAND_144[6:0];
  _RAND_145 = {1{`RANDOM}};
  rob_uop_8_stale_dst = _RAND_145[6:0];
  _RAND_146 = {1{`RANDOM}};
  rob_uop_8_arch_dst = _RAND_146[4:0];
  _RAND_147 = {2{`RANDOM}};
  rob_uop_8_dst_value = _RAND_147[63:0];
  _RAND_148 = {2{`RANDOM}};
  rob_uop_8_src1_value = _RAND_148[63:0];
  _RAND_149 = {1{`RANDOM}};
  rob_uop_8_alu_sel = _RAND_149[4:0];
  _RAND_150 = {1{`RANDOM}};
  rob_uop_9_pc = _RAND_150[31:0];
  _RAND_151 = {1{`RANDOM}};
  rob_uop_9_inst = _RAND_151[31:0];
  _RAND_152 = {1{`RANDOM}};
  rob_uop_9_func_code = _RAND_152[6:0];
  _RAND_153 = {1{`RANDOM}};
  rob_uop_9_phy_dst = _RAND_153[6:0];
  _RAND_154 = {1{`RANDOM}};
  rob_uop_9_stale_dst = _RAND_154[6:0];
  _RAND_155 = {1{`RANDOM}};
  rob_uop_9_arch_dst = _RAND_155[4:0];
  _RAND_156 = {2{`RANDOM}};
  rob_uop_9_dst_value = _RAND_156[63:0];
  _RAND_157 = {2{`RANDOM}};
  rob_uop_9_src1_value = _RAND_157[63:0];
  _RAND_158 = {1{`RANDOM}};
  rob_uop_9_alu_sel = _RAND_158[4:0];
  _RAND_159 = {1{`RANDOM}};
  rob_uop_10_pc = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  rob_uop_10_inst = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  rob_uop_10_func_code = _RAND_161[6:0];
  _RAND_162 = {1{`RANDOM}};
  rob_uop_10_phy_dst = _RAND_162[6:0];
  _RAND_163 = {1{`RANDOM}};
  rob_uop_10_stale_dst = _RAND_163[6:0];
  _RAND_164 = {1{`RANDOM}};
  rob_uop_10_arch_dst = _RAND_164[4:0];
  _RAND_165 = {2{`RANDOM}};
  rob_uop_10_dst_value = _RAND_165[63:0];
  _RAND_166 = {2{`RANDOM}};
  rob_uop_10_src1_value = _RAND_166[63:0];
  _RAND_167 = {1{`RANDOM}};
  rob_uop_10_alu_sel = _RAND_167[4:0];
  _RAND_168 = {1{`RANDOM}};
  rob_uop_11_pc = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  rob_uop_11_inst = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  rob_uop_11_func_code = _RAND_170[6:0];
  _RAND_171 = {1{`RANDOM}};
  rob_uop_11_phy_dst = _RAND_171[6:0];
  _RAND_172 = {1{`RANDOM}};
  rob_uop_11_stale_dst = _RAND_172[6:0];
  _RAND_173 = {1{`RANDOM}};
  rob_uop_11_arch_dst = _RAND_173[4:0];
  _RAND_174 = {2{`RANDOM}};
  rob_uop_11_dst_value = _RAND_174[63:0];
  _RAND_175 = {2{`RANDOM}};
  rob_uop_11_src1_value = _RAND_175[63:0];
  _RAND_176 = {1{`RANDOM}};
  rob_uop_11_alu_sel = _RAND_176[4:0];
  _RAND_177 = {1{`RANDOM}};
  rob_uop_12_pc = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  rob_uop_12_inst = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  rob_uop_12_func_code = _RAND_179[6:0];
  _RAND_180 = {1{`RANDOM}};
  rob_uop_12_phy_dst = _RAND_180[6:0];
  _RAND_181 = {1{`RANDOM}};
  rob_uop_12_stale_dst = _RAND_181[6:0];
  _RAND_182 = {1{`RANDOM}};
  rob_uop_12_arch_dst = _RAND_182[4:0];
  _RAND_183 = {2{`RANDOM}};
  rob_uop_12_dst_value = _RAND_183[63:0];
  _RAND_184 = {2{`RANDOM}};
  rob_uop_12_src1_value = _RAND_184[63:0];
  _RAND_185 = {1{`RANDOM}};
  rob_uop_12_alu_sel = _RAND_185[4:0];
  _RAND_186 = {1{`RANDOM}};
  rob_uop_13_pc = _RAND_186[31:0];
  _RAND_187 = {1{`RANDOM}};
  rob_uop_13_inst = _RAND_187[31:0];
  _RAND_188 = {1{`RANDOM}};
  rob_uop_13_func_code = _RAND_188[6:0];
  _RAND_189 = {1{`RANDOM}};
  rob_uop_13_phy_dst = _RAND_189[6:0];
  _RAND_190 = {1{`RANDOM}};
  rob_uop_13_stale_dst = _RAND_190[6:0];
  _RAND_191 = {1{`RANDOM}};
  rob_uop_13_arch_dst = _RAND_191[4:0];
  _RAND_192 = {2{`RANDOM}};
  rob_uop_13_dst_value = _RAND_192[63:0];
  _RAND_193 = {2{`RANDOM}};
  rob_uop_13_src1_value = _RAND_193[63:0];
  _RAND_194 = {1{`RANDOM}};
  rob_uop_13_alu_sel = _RAND_194[4:0];
  _RAND_195 = {1{`RANDOM}};
  rob_uop_14_pc = _RAND_195[31:0];
  _RAND_196 = {1{`RANDOM}};
  rob_uop_14_inst = _RAND_196[31:0];
  _RAND_197 = {1{`RANDOM}};
  rob_uop_14_func_code = _RAND_197[6:0];
  _RAND_198 = {1{`RANDOM}};
  rob_uop_14_phy_dst = _RAND_198[6:0];
  _RAND_199 = {1{`RANDOM}};
  rob_uop_14_stale_dst = _RAND_199[6:0];
  _RAND_200 = {1{`RANDOM}};
  rob_uop_14_arch_dst = _RAND_200[4:0];
  _RAND_201 = {2{`RANDOM}};
  rob_uop_14_dst_value = _RAND_201[63:0];
  _RAND_202 = {2{`RANDOM}};
  rob_uop_14_src1_value = _RAND_202[63:0];
  _RAND_203 = {1{`RANDOM}};
  rob_uop_14_alu_sel = _RAND_203[4:0];
  _RAND_204 = {1{`RANDOM}};
  rob_uop_15_pc = _RAND_204[31:0];
  _RAND_205 = {1{`RANDOM}};
  rob_uop_15_inst = _RAND_205[31:0];
  _RAND_206 = {1{`RANDOM}};
  rob_uop_15_func_code = _RAND_206[6:0];
  _RAND_207 = {1{`RANDOM}};
  rob_uop_15_phy_dst = _RAND_207[6:0];
  _RAND_208 = {1{`RANDOM}};
  rob_uop_15_stale_dst = _RAND_208[6:0];
  _RAND_209 = {1{`RANDOM}};
  rob_uop_15_arch_dst = _RAND_209[4:0];
  _RAND_210 = {2{`RANDOM}};
  rob_uop_15_dst_value = _RAND_210[63:0];
  _RAND_211 = {2{`RANDOM}};
  rob_uop_15_src1_value = _RAND_211[63:0];
  _RAND_212 = {1{`RANDOM}};
  rob_uop_15_alu_sel = _RAND_212[4:0];
  _RAND_213 = {1{`RANDOM}};
  rob_uop_16_pc = _RAND_213[31:0];
  _RAND_214 = {1{`RANDOM}};
  rob_uop_16_inst = _RAND_214[31:0];
  _RAND_215 = {1{`RANDOM}};
  rob_uop_16_func_code = _RAND_215[6:0];
  _RAND_216 = {1{`RANDOM}};
  rob_uop_16_phy_dst = _RAND_216[6:0];
  _RAND_217 = {1{`RANDOM}};
  rob_uop_16_stale_dst = _RAND_217[6:0];
  _RAND_218 = {1{`RANDOM}};
  rob_uop_16_arch_dst = _RAND_218[4:0];
  _RAND_219 = {2{`RANDOM}};
  rob_uop_16_dst_value = _RAND_219[63:0];
  _RAND_220 = {2{`RANDOM}};
  rob_uop_16_src1_value = _RAND_220[63:0];
  _RAND_221 = {1{`RANDOM}};
  rob_uop_16_alu_sel = _RAND_221[4:0];
  _RAND_222 = {1{`RANDOM}};
  rob_uop_17_pc = _RAND_222[31:0];
  _RAND_223 = {1{`RANDOM}};
  rob_uop_17_inst = _RAND_223[31:0];
  _RAND_224 = {1{`RANDOM}};
  rob_uop_17_func_code = _RAND_224[6:0];
  _RAND_225 = {1{`RANDOM}};
  rob_uop_17_phy_dst = _RAND_225[6:0];
  _RAND_226 = {1{`RANDOM}};
  rob_uop_17_stale_dst = _RAND_226[6:0];
  _RAND_227 = {1{`RANDOM}};
  rob_uop_17_arch_dst = _RAND_227[4:0];
  _RAND_228 = {2{`RANDOM}};
  rob_uop_17_dst_value = _RAND_228[63:0];
  _RAND_229 = {2{`RANDOM}};
  rob_uop_17_src1_value = _RAND_229[63:0];
  _RAND_230 = {1{`RANDOM}};
  rob_uop_17_alu_sel = _RAND_230[4:0];
  _RAND_231 = {1{`RANDOM}};
  rob_uop_18_pc = _RAND_231[31:0];
  _RAND_232 = {1{`RANDOM}};
  rob_uop_18_inst = _RAND_232[31:0];
  _RAND_233 = {1{`RANDOM}};
  rob_uop_18_func_code = _RAND_233[6:0];
  _RAND_234 = {1{`RANDOM}};
  rob_uop_18_phy_dst = _RAND_234[6:0];
  _RAND_235 = {1{`RANDOM}};
  rob_uop_18_stale_dst = _RAND_235[6:0];
  _RAND_236 = {1{`RANDOM}};
  rob_uop_18_arch_dst = _RAND_236[4:0];
  _RAND_237 = {2{`RANDOM}};
  rob_uop_18_dst_value = _RAND_237[63:0];
  _RAND_238 = {2{`RANDOM}};
  rob_uop_18_src1_value = _RAND_238[63:0];
  _RAND_239 = {1{`RANDOM}};
  rob_uop_18_alu_sel = _RAND_239[4:0];
  _RAND_240 = {1{`RANDOM}};
  rob_uop_19_pc = _RAND_240[31:0];
  _RAND_241 = {1{`RANDOM}};
  rob_uop_19_inst = _RAND_241[31:0];
  _RAND_242 = {1{`RANDOM}};
  rob_uop_19_func_code = _RAND_242[6:0];
  _RAND_243 = {1{`RANDOM}};
  rob_uop_19_phy_dst = _RAND_243[6:0];
  _RAND_244 = {1{`RANDOM}};
  rob_uop_19_stale_dst = _RAND_244[6:0];
  _RAND_245 = {1{`RANDOM}};
  rob_uop_19_arch_dst = _RAND_245[4:0];
  _RAND_246 = {2{`RANDOM}};
  rob_uop_19_dst_value = _RAND_246[63:0];
  _RAND_247 = {2{`RANDOM}};
  rob_uop_19_src1_value = _RAND_247[63:0];
  _RAND_248 = {1{`RANDOM}};
  rob_uop_19_alu_sel = _RAND_248[4:0];
  _RAND_249 = {1{`RANDOM}};
  rob_uop_20_pc = _RAND_249[31:0];
  _RAND_250 = {1{`RANDOM}};
  rob_uop_20_inst = _RAND_250[31:0];
  _RAND_251 = {1{`RANDOM}};
  rob_uop_20_func_code = _RAND_251[6:0];
  _RAND_252 = {1{`RANDOM}};
  rob_uop_20_phy_dst = _RAND_252[6:0];
  _RAND_253 = {1{`RANDOM}};
  rob_uop_20_stale_dst = _RAND_253[6:0];
  _RAND_254 = {1{`RANDOM}};
  rob_uop_20_arch_dst = _RAND_254[4:0];
  _RAND_255 = {2{`RANDOM}};
  rob_uop_20_dst_value = _RAND_255[63:0];
  _RAND_256 = {2{`RANDOM}};
  rob_uop_20_src1_value = _RAND_256[63:0];
  _RAND_257 = {1{`RANDOM}};
  rob_uop_20_alu_sel = _RAND_257[4:0];
  _RAND_258 = {1{`RANDOM}};
  rob_uop_21_pc = _RAND_258[31:0];
  _RAND_259 = {1{`RANDOM}};
  rob_uop_21_inst = _RAND_259[31:0];
  _RAND_260 = {1{`RANDOM}};
  rob_uop_21_func_code = _RAND_260[6:0];
  _RAND_261 = {1{`RANDOM}};
  rob_uop_21_phy_dst = _RAND_261[6:0];
  _RAND_262 = {1{`RANDOM}};
  rob_uop_21_stale_dst = _RAND_262[6:0];
  _RAND_263 = {1{`RANDOM}};
  rob_uop_21_arch_dst = _RAND_263[4:0];
  _RAND_264 = {2{`RANDOM}};
  rob_uop_21_dst_value = _RAND_264[63:0];
  _RAND_265 = {2{`RANDOM}};
  rob_uop_21_src1_value = _RAND_265[63:0];
  _RAND_266 = {1{`RANDOM}};
  rob_uop_21_alu_sel = _RAND_266[4:0];
  _RAND_267 = {1{`RANDOM}};
  rob_uop_22_pc = _RAND_267[31:0];
  _RAND_268 = {1{`RANDOM}};
  rob_uop_22_inst = _RAND_268[31:0];
  _RAND_269 = {1{`RANDOM}};
  rob_uop_22_func_code = _RAND_269[6:0];
  _RAND_270 = {1{`RANDOM}};
  rob_uop_22_phy_dst = _RAND_270[6:0];
  _RAND_271 = {1{`RANDOM}};
  rob_uop_22_stale_dst = _RAND_271[6:0];
  _RAND_272 = {1{`RANDOM}};
  rob_uop_22_arch_dst = _RAND_272[4:0];
  _RAND_273 = {2{`RANDOM}};
  rob_uop_22_dst_value = _RAND_273[63:0];
  _RAND_274 = {2{`RANDOM}};
  rob_uop_22_src1_value = _RAND_274[63:0];
  _RAND_275 = {1{`RANDOM}};
  rob_uop_22_alu_sel = _RAND_275[4:0];
  _RAND_276 = {1{`RANDOM}};
  rob_uop_23_pc = _RAND_276[31:0];
  _RAND_277 = {1{`RANDOM}};
  rob_uop_23_inst = _RAND_277[31:0];
  _RAND_278 = {1{`RANDOM}};
  rob_uop_23_func_code = _RAND_278[6:0];
  _RAND_279 = {1{`RANDOM}};
  rob_uop_23_phy_dst = _RAND_279[6:0];
  _RAND_280 = {1{`RANDOM}};
  rob_uop_23_stale_dst = _RAND_280[6:0];
  _RAND_281 = {1{`RANDOM}};
  rob_uop_23_arch_dst = _RAND_281[4:0];
  _RAND_282 = {2{`RANDOM}};
  rob_uop_23_dst_value = _RAND_282[63:0];
  _RAND_283 = {2{`RANDOM}};
  rob_uop_23_src1_value = _RAND_283[63:0];
  _RAND_284 = {1{`RANDOM}};
  rob_uop_23_alu_sel = _RAND_284[4:0];
  _RAND_285 = {1{`RANDOM}};
  rob_uop_24_pc = _RAND_285[31:0];
  _RAND_286 = {1{`RANDOM}};
  rob_uop_24_inst = _RAND_286[31:0];
  _RAND_287 = {1{`RANDOM}};
  rob_uop_24_func_code = _RAND_287[6:0];
  _RAND_288 = {1{`RANDOM}};
  rob_uop_24_phy_dst = _RAND_288[6:0];
  _RAND_289 = {1{`RANDOM}};
  rob_uop_24_stale_dst = _RAND_289[6:0];
  _RAND_290 = {1{`RANDOM}};
  rob_uop_24_arch_dst = _RAND_290[4:0];
  _RAND_291 = {2{`RANDOM}};
  rob_uop_24_dst_value = _RAND_291[63:0];
  _RAND_292 = {2{`RANDOM}};
  rob_uop_24_src1_value = _RAND_292[63:0];
  _RAND_293 = {1{`RANDOM}};
  rob_uop_24_alu_sel = _RAND_293[4:0];
  _RAND_294 = {1{`RANDOM}};
  rob_uop_25_pc = _RAND_294[31:0];
  _RAND_295 = {1{`RANDOM}};
  rob_uop_25_inst = _RAND_295[31:0];
  _RAND_296 = {1{`RANDOM}};
  rob_uop_25_func_code = _RAND_296[6:0];
  _RAND_297 = {1{`RANDOM}};
  rob_uop_25_phy_dst = _RAND_297[6:0];
  _RAND_298 = {1{`RANDOM}};
  rob_uop_25_stale_dst = _RAND_298[6:0];
  _RAND_299 = {1{`RANDOM}};
  rob_uop_25_arch_dst = _RAND_299[4:0];
  _RAND_300 = {2{`RANDOM}};
  rob_uop_25_dst_value = _RAND_300[63:0];
  _RAND_301 = {2{`RANDOM}};
  rob_uop_25_src1_value = _RAND_301[63:0];
  _RAND_302 = {1{`RANDOM}};
  rob_uop_25_alu_sel = _RAND_302[4:0];
  _RAND_303 = {1{`RANDOM}};
  rob_uop_26_pc = _RAND_303[31:0];
  _RAND_304 = {1{`RANDOM}};
  rob_uop_26_inst = _RAND_304[31:0];
  _RAND_305 = {1{`RANDOM}};
  rob_uop_26_func_code = _RAND_305[6:0];
  _RAND_306 = {1{`RANDOM}};
  rob_uop_26_phy_dst = _RAND_306[6:0];
  _RAND_307 = {1{`RANDOM}};
  rob_uop_26_stale_dst = _RAND_307[6:0];
  _RAND_308 = {1{`RANDOM}};
  rob_uop_26_arch_dst = _RAND_308[4:0];
  _RAND_309 = {2{`RANDOM}};
  rob_uop_26_dst_value = _RAND_309[63:0];
  _RAND_310 = {2{`RANDOM}};
  rob_uop_26_src1_value = _RAND_310[63:0];
  _RAND_311 = {1{`RANDOM}};
  rob_uop_26_alu_sel = _RAND_311[4:0];
  _RAND_312 = {1{`RANDOM}};
  rob_uop_27_pc = _RAND_312[31:0];
  _RAND_313 = {1{`RANDOM}};
  rob_uop_27_inst = _RAND_313[31:0];
  _RAND_314 = {1{`RANDOM}};
  rob_uop_27_func_code = _RAND_314[6:0];
  _RAND_315 = {1{`RANDOM}};
  rob_uop_27_phy_dst = _RAND_315[6:0];
  _RAND_316 = {1{`RANDOM}};
  rob_uop_27_stale_dst = _RAND_316[6:0];
  _RAND_317 = {1{`RANDOM}};
  rob_uop_27_arch_dst = _RAND_317[4:0];
  _RAND_318 = {2{`RANDOM}};
  rob_uop_27_dst_value = _RAND_318[63:0];
  _RAND_319 = {2{`RANDOM}};
  rob_uop_27_src1_value = _RAND_319[63:0];
  _RAND_320 = {1{`RANDOM}};
  rob_uop_27_alu_sel = _RAND_320[4:0];
  _RAND_321 = {1{`RANDOM}};
  rob_uop_28_pc = _RAND_321[31:0];
  _RAND_322 = {1{`RANDOM}};
  rob_uop_28_inst = _RAND_322[31:0];
  _RAND_323 = {1{`RANDOM}};
  rob_uop_28_func_code = _RAND_323[6:0];
  _RAND_324 = {1{`RANDOM}};
  rob_uop_28_phy_dst = _RAND_324[6:0];
  _RAND_325 = {1{`RANDOM}};
  rob_uop_28_stale_dst = _RAND_325[6:0];
  _RAND_326 = {1{`RANDOM}};
  rob_uop_28_arch_dst = _RAND_326[4:0];
  _RAND_327 = {2{`RANDOM}};
  rob_uop_28_dst_value = _RAND_327[63:0];
  _RAND_328 = {2{`RANDOM}};
  rob_uop_28_src1_value = _RAND_328[63:0];
  _RAND_329 = {1{`RANDOM}};
  rob_uop_28_alu_sel = _RAND_329[4:0];
  _RAND_330 = {1{`RANDOM}};
  rob_uop_29_pc = _RAND_330[31:0];
  _RAND_331 = {1{`RANDOM}};
  rob_uop_29_inst = _RAND_331[31:0];
  _RAND_332 = {1{`RANDOM}};
  rob_uop_29_func_code = _RAND_332[6:0];
  _RAND_333 = {1{`RANDOM}};
  rob_uop_29_phy_dst = _RAND_333[6:0];
  _RAND_334 = {1{`RANDOM}};
  rob_uop_29_stale_dst = _RAND_334[6:0];
  _RAND_335 = {1{`RANDOM}};
  rob_uop_29_arch_dst = _RAND_335[4:0];
  _RAND_336 = {2{`RANDOM}};
  rob_uop_29_dst_value = _RAND_336[63:0];
  _RAND_337 = {2{`RANDOM}};
  rob_uop_29_src1_value = _RAND_337[63:0];
  _RAND_338 = {1{`RANDOM}};
  rob_uop_29_alu_sel = _RAND_338[4:0];
  _RAND_339 = {1{`RANDOM}};
  rob_uop_30_pc = _RAND_339[31:0];
  _RAND_340 = {1{`RANDOM}};
  rob_uop_30_inst = _RAND_340[31:0];
  _RAND_341 = {1{`RANDOM}};
  rob_uop_30_func_code = _RAND_341[6:0];
  _RAND_342 = {1{`RANDOM}};
  rob_uop_30_phy_dst = _RAND_342[6:0];
  _RAND_343 = {1{`RANDOM}};
  rob_uop_30_stale_dst = _RAND_343[6:0];
  _RAND_344 = {1{`RANDOM}};
  rob_uop_30_arch_dst = _RAND_344[4:0];
  _RAND_345 = {2{`RANDOM}};
  rob_uop_30_dst_value = _RAND_345[63:0];
  _RAND_346 = {2{`RANDOM}};
  rob_uop_30_src1_value = _RAND_346[63:0];
  _RAND_347 = {1{`RANDOM}};
  rob_uop_30_alu_sel = _RAND_347[4:0];
  _RAND_348 = {1{`RANDOM}};
  rob_uop_31_pc = _RAND_348[31:0];
  _RAND_349 = {1{`RANDOM}};
  rob_uop_31_inst = _RAND_349[31:0];
  _RAND_350 = {1{`RANDOM}};
  rob_uop_31_func_code = _RAND_350[6:0];
  _RAND_351 = {1{`RANDOM}};
  rob_uop_31_phy_dst = _RAND_351[6:0];
  _RAND_352 = {1{`RANDOM}};
  rob_uop_31_stale_dst = _RAND_352[6:0];
  _RAND_353 = {1{`RANDOM}};
  rob_uop_31_arch_dst = _RAND_353[4:0];
  _RAND_354 = {2{`RANDOM}};
  rob_uop_31_dst_value = _RAND_354[63:0];
  _RAND_355 = {2{`RANDOM}};
  rob_uop_31_src1_value = _RAND_355[63:0];
  _RAND_356 = {1{`RANDOM}};
  rob_uop_31_alu_sel = _RAND_356[4:0];
  _RAND_357 = {1{`RANDOM}};
  rob_uop_32_pc = _RAND_357[31:0];
  _RAND_358 = {1{`RANDOM}};
  rob_uop_32_inst = _RAND_358[31:0];
  _RAND_359 = {1{`RANDOM}};
  rob_uop_32_func_code = _RAND_359[6:0];
  _RAND_360 = {1{`RANDOM}};
  rob_uop_32_phy_dst = _RAND_360[6:0];
  _RAND_361 = {1{`RANDOM}};
  rob_uop_32_stale_dst = _RAND_361[6:0];
  _RAND_362 = {1{`RANDOM}};
  rob_uop_32_arch_dst = _RAND_362[4:0];
  _RAND_363 = {2{`RANDOM}};
  rob_uop_32_dst_value = _RAND_363[63:0];
  _RAND_364 = {2{`RANDOM}};
  rob_uop_32_src1_value = _RAND_364[63:0];
  _RAND_365 = {1{`RANDOM}};
  rob_uop_32_alu_sel = _RAND_365[4:0];
  _RAND_366 = {1{`RANDOM}};
  rob_uop_33_pc = _RAND_366[31:0];
  _RAND_367 = {1{`RANDOM}};
  rob_uop_33_inst = _RAND_367[31:0];
  _RAND_368 = {1{`RANDOM}};
  rob_uop_33_func_code = _RAND_368[6:0];
  _RAND_369 = {1{`RANDOM}};
  rob_uop_33_phy_dst = _RAND_369[6:0];
  _RAND_370 = {1{`RANDOM}};
  rob_uop_33_stale_dst = _RAND_370[6:0];
  _RAND_371 = {1{`RANDOM}};
  rob_uop_33_arch_dst = _RAND_371[4:0];
  _RAND_372 = {2{`RANDOM}};
  rob_uop_33_dst_value = _RAND_372[63:0];
  _RAND_373 = {2{`RANDOM}};
  rob_uop_33_src1_value = _RAND_373[63:0];
  _RAND_374 = {1{`RANDOM}};
  rob_uop_33_alu_sel = _RAND_374[4:0];
  _RAND_375 = {1{`RANDOM}};
  rob_uop_34_pc = _RAND_375[31:0];
  _RAND_376 = {1{`RANDOM}};
  rob_uop_34_inst = _RAND_376[31:0];
  _RAND_377 = {1{`RANDOM}};
  rob_uop_34_func_code = _RAND_377[6:0];
  _RAND_378 = {1{`RANDOM}};
  rob_uop_34_phy_dst = _RAND_378[6:0];
  _RAND_379 = {1{`RANDOM}};
  rob_uop_34_stale_dst = _RAND_379[6:0];
  _RAND_380 = {1{`RANDOM}};
  rob_uop_34_arch_dst = _RAND_380[4:0];
  _RAND_381 = {2{`RANDOM}};
  rob_uop_34_dst_value = _RAND_381[63:0];
  _RAND_382 = {2{`RANDOM}};
  rob_uop_34_src1_value = _RAND_382[63:0];
  _RAND_383 = {1{`RANDOM}};
  rob_uop_34_alu_sel = _RAND_383[4:0];
  _RAND_384 = {1{`RANDOM}};
  rob_uop_35_pc = _RAND_384[31:0];
  _RAND_385 = {1{`RANDOM}};
  rob_uop_35_inst = _RAND_385[31:0];
  _RAND_386 = {1{`RANDOM}};
  rob_uop_35_func_code = _RAND_386[6:0];
  _RAND_387 = {1{`RANDOM}};
  rob_uop_35_phy_dst = _RAND_387[6:0];
  _RAND_388 = {1{`RANDOM}};
  rob_uop_35_stale_dst = _RAND_388[6:0];
  _RAND_389 = {1{`RANDOM}};
  rob_uop_35_arch_dst = _RAND_389[4:0];
  _RAND_390 = {2{`RANDOM}};
  rob_uop_35_dst_value = _RAND_390[63:0];
  _RAND_391 = {2{`RANDOM}};
  rob_uop_35_src1_value = _RAND_391[63:0];
  _RAND_392 = {1{`RANDOM}};
  rob_uop_35_alu_sel = _RAND_392[4:0];
  _RAND_393 = {1{`RANDOM}};
  rob_uop_36_pc = _RAND_393[31:0];
  _RAND_394 = {1{`RANDOM}};
  rob_uop_36_inst = _RAND_394[31:0];
  _RAND_395 = {1{`RANDOM}};
  rob_uop_36_func_code = _RAND_395[6:0];
  _RAND_396 = {1{`RANDOM}};
  rob_uop_36_phy_dst = _RAND_396[6:0];
  _RAND_397 = {1{`RANDOM}};
  rob_uop_36_stale_dst = _RAND_397[6:0];
  _RAND_398 = {1{`RANDOM}};
  rob_uop_36_arch_dst = _RAND_398[4:0];
  _RAND_399 = {2{`RANDOM}};
  rob_uop_36_dst_value = _RAND_399[63:0];
  _RAND_400 = {2{`RANDOM}};
  rob_uop_36_src1_value = _RAND_400[63:0];
  _RAND_401 = {1{`RANDOM}};
  rob_uop_36_alu_sel = _RAND_401[4:0];
  _RAND_402 = {1{`RANDOM}};
  rob_uop_37_pc = _RAND_402[31:0];
  _RAND_403 = {1{`RANDOM}};
  rob_uop_37_inst = _RAND_403[31:0];
  _RAND_404 = {1{`RANDOM}};
  rob_uop_37_func_code = _RAND_404[6:0];
  _RAND_405 = {1{`RANDOM}};
  rob_uop_37_phy_dst = _RAND_405[6:0];
  _RAND_406 = {1{`RANDOM}};
  rob_uop_37_stale_dst = _RAND_406[6:0];
  _RAND_407 = {1{`RANDOM}};
  rob_uop_37_arch_dst = _RAND_407[4:0];
  _RAND_408 = {2{`RANDOM}};
  rob_uop_37_dst_value = _RAND_408[63:0];
  _RAND_409 = {2{`RANDOM}};
  rob_uop_37_src1_value = _RAND_409[63:0];
  _RAND_410 = {1{`RANDOM}};
  rob_uop_37_alu_sel = _RAND_410[4:0];
  _RAND_411 = {1{`RANDOM}};
  rob_uop_38_pc = _RAND_411[31:0];
  _RAND_412 = {1{`RANDOM}};
  rob_uop_38_inst = _RAND_412[31:0];
  _RAND_413 = {1{`RANDOM}};
  rob_uop_38_func_code = _RAND_413[6:0];
  _RAND_414 = {1{`RANDOM}};
  rob_uop_38_phy_dst = _RAND_414[6:0];
  _RAND_415 = {1{`RANDOM}};
  rob_uop_38_stale_dst = _RAND_415[6:0];
  _RAND_416 = {1{`RANDOM}};
  rob_uop_38_arch_dst = _RAND_416[4:0];
  _RAND_417 = {2{`RANDOM}};
  rob_uop_38_dst_value = _RAND_417[63:0];
  _RAND_418 = {2{`RANDOM}};
  rob_uop_38_src1_value = _RAND_418[63:0];
  _RAND_419 = {1{`RANDOM}};
  rob_uop_38_alu_sel = _RAND_419[4:0];
  _RAND_420 = {1{`RANDOM}};
  rob_uop_39_pc = _RAND_420[31:0];
  _RAND_421 = {1{`RANDOM}};
  rob_uop_39_inst = _RAND_421[31:0];
  _RAND_422 = {1{`RANDOM}};
  rob_uop_39_func_code = _RAND_422[6:0];
  _RAND_423 = {1{`RANDOM}};
  rob_uop_39_phy_dst = _RAND_423[6:0];
  _RAND_424 = {1{`RANDOM}};
  rob_uop_39_stale_dst = _RAND_424[6:0];
  _RAND_425 = {1{`RANDOM}};
  rob_uop_39_arch_dst = _RAND_425[4:0];
  _RAND_426 = {2{`RANDOM}};
  rob_uop_39_dst_value = _RAND_426[63:0];
  _RAND_427 = {2{`RANDOM}};
  rob_uop_39_src1_value = _RAND_427[63:0];
  _RAND_428 = {1{`RANDOM}};
  rob_uop_39_alu_sel = _RAND_428[4:0];
  _RAND_429 = {1{`RANDOM}};
  rob_uop_40_pc = _RAND_429[31:0];
  _RAND_430 = {1{`RANDOM}};
  rob_uop_40_inst = _RAND_430[31:0];
  _RAND_431 = {1{`RANDOM}};
  rob_uop_40_func_code = _RAND_431[6:0];
  _RAND_432 = {1{`RANDOM}};
  rob_uop_40_phy_dst = _RAND_432[6:0];
  _RAND_433 = {1{`RANDOM}};
  rob_uop_40_stale_dst = _RAND_433[6:0];
  _RAND_434 = {1{`RANDOM}};
  rob_uop_40_arch_dst = _RAND_434[4:0];
  _RAND_435 = {2{`RANDOM}};
  rob_uop_40_dst_value = _RAND_435[63:0];
  _RAND_436 = {2{`RANDOM}};
  rob_uop_40_src1_value = _RAND_436[63:0];
  _RAND_437 = {1{`RANDOM}};
  rob_uop_40_alu_sel = _RAND_437[4:0];
  _RAND_438 = {1{`RANDOM}};
  rob_uop_41_pc = _RAND_438[31:0];
  _RAND_439 = {1{`RANDOM}};
  rob_uop_41_inst = _RAND_439[31:0];
  _RAND_440 = {1{`RANDOM}};
  rob_uop_41_func_code = _RAND_440[6:0];
  _RAND_441 = {1{`RANDOM}};
  rob_uop_41_phy_dst = _RAND_441[6:0];
  _RAND_442 = {1{`RANDOM}};
  rob_uop_41_stale_dst = _RAND_442[6:0];
  _RAND_443 = {1{`RANDOM}};
  rob_uop_41_arch_dst = _RAND_443[4:0];
  _RAND_444 = {2{`RANDOM}};
  rob_uop_41_dst_value = _RAND_444[63:0];
  _RAND_445 = {2{`RANDOM}};
  rob_uop_41_src1_value = _RAND_445[63:0];
  _RAND_446 = {1{`RANDOM}};
  rob_uop_41_alu_sel = _RAND_446[4:0];
  _RAND_447 = {1{`RANDOM}};
  rob_uop_42_pc = _RAND_447[31:0];
  _RAND_448 = {1{`RANDOM}};
  rob_uop_42_inst = _RAND_448[31:0];
  _RAND_449 = {1{`RANDOM}};
  rob_uop_42_func_code = _RAND_449[6:0];
  _RAND_450 = {1{`RANDOM}};
  rob_uop_42_phy_dst = _RAND_450[6:0];
  _RAND_451 = {1{`RANDOM}};
  rob_uop_42_stale_dst = _RAND_451[6:0];
  _RAND_452 = {1{`RANDOM}};
  rob_uop_42_arch_dst = _RAND_452[4:0];
  _RAND_453 = {2{`RANDOM}};
  rob_uop_42_dst_value = _RAND_453[63:0];
  _RAND_454 = {2{`RANDOM}};
  rob_uop_42_src1_value = _RAND_454[63:0];
  _RAND_455 = {1{`RANDOM}};
  rob_uop_42_alu_sel = _RAND_455[4:0];
  _RAND_456 = {1{`RANDOM}};
  rob_uop_43_pc = _RAND_456[31:0];
  _RAND_457 = {1{`RANDOM}};
  rob_uop_43_inst = _RAND_457[31:0];
  _RAND_458 = {1{`RANDOM}};
  rob_uop_43_func_code = _RAND_458[6:0];
  _RAND_459 = {1{`RANDOM}};
  rob_uop_43_phy_dst = _RAND_459[6:0];
  _RAND_460 = {1{`RANDOM}};
  rob_uop_43_stale_dst = _RAND_460[6:0];
  _RAND_461 = {1{`RANDOM}};
  rob_uop_43_arch_dst = _RAND_461[4:0];
  _RAND_462 = {2{`RANDOM}};
  rob_uop_43_dst_value = _RAND_462[63:0];
  _RAND_463 = {2{`RANDOM}};
  rob_uop_43_src1_value = _RAND_463[63:0];
  _RAND_464 = {1{`RANDOM}};
  rob_uop_43_alu_sel = _RAND_464[4:0];
  _RAND_465 = {1{`RANDOM}};
  rob_uop_44_pc = _RAND_465[31:0];
  _RAND_466 = {1{`RANDOM}};
  rob_uop_44_inst = _RAND_466[31:0];
  _RAND_467 = {1{`RANDOM}};
  rob_uop_44_func_code = _RAND_467[6:0];
  _RAND_468 = {1{`RANDOM}};
  rob_uop_44_phy_dst = _RAND_468[6:0];
  _RAND_469 = {1{`RANDOM}};
  rob_uop_44_stale_dst = _RAND_469[6:0];
  _RAND_470 = {1{`RANDOM}};
  rob_uop_44_arch_dst = _RAND_470[4:0];
  _RAND_471 = {2{`RANDOM}};
  rob_uop_44_dst_value = _RAND_471[63:0];
  _RAND_472 = {2{`RANDOM}};
  rob_uop_44_src1_value = _RAND_472[63:0];
  _RAND_473 = {1{`RANDOM}};
  rob_uop_44_alu_sel = _RAND_473[4:0];
  _RAND_474 = {1{`RANDOM}};
  rob_uop_45_pc = _RAND_474[31:0];
  _RAND_475 = {1{`RANDOM}};
  rob_uop_45_inst = _RAND_475[31:0];
  _RAND_476 = {1{`RANDOM}};
  rob_uop_45_func_code = _RAND_476[6:0];
  _RAND_477 = {1{`RANDOM}};
  rob_uop_45_phy_dst = _RAND_477[6:0];
  _RAND_478 = {1{`RANDOM}};
  rob_uop_45_stale_dst = _RAND_478[6:0];
  _RAND_479 = {1{`RANDOM}};
  rob_uop_45_arch_dst = _RAND_479[4:0];
  _RAND_480 = {2{`RANDOM}};
  rob_uop_45_dst_value = _RAND_480[63:0];
  _RAND_481 = {2{`RANDOM}};
  rob_uop_45_src1_value = _RAND_481[63:0];
  _RAND_482 = {1{`RANDOM}};
  rob_uop_45_alu_sel = _RAND_482[4:0];
  _RAND_483 = {1{`RANDOM}};
  rob_uop_46_pc = _RAND_483[31:0];
  _RAND_484 = {1{`RANDOM}};
  rob_uop_46_inst = _RAND_484[31:0];
  _RAND_485 = {1{`RANDOM}};
  rob_uop_46_func_code = _RAND_485[6:0];
  _RAND_486 = {1{`RANDOM}};
  rob_uop_46_phy_dst = _RAND_486[6:0];
  _RAND_487 = {1{`RANDOM}};
  rob_uop_46_stale_dst = _RAND_487[6:0];
  _RAND_488 = {1{`RANDOM}};
  rob_uop_46_arch_dst = _RAND_488[4:0];
  _RAND_489 = {2{`RANDOM}};
  rob_uop_46_dst_value = _RAND_489[63:0];
  _RAND_490 = {2{`RANDOM}};
  rob_uop_46_src1_value = _RAND_490[63:0];
  _RAND_491 = {1{`RANDOM}};
  rob_uop_46_alu_sel = _RAND_491[4:0];
  _RAND_492 = {1{`RANDOM}};
  rob_uop_47_pc = _RAND_492[31:0];
  _RAND_493 = {1{`RANDOM}};
  rob_uop_47_inst = _RAND_493[31:0];
  _RAND_494 = {1{`RANDOM}};
  rob_uop_47_func_code = _RAND_494[6:0];
  _RAND_495 = {1{`RANDOM}};
  rob_uop_47_phy_dst = _RAND_495[6:0];
  _RAND_496 = {1{`RANDOM}};
  rob_uop_47_stale_dst = _RAND_496[6:0];
  _RAND_497 = {1{`RANDOM}};
  rob_uop_47_arch_dst = _RAND_497[4:0];
  _RAND_498 = {2{`RANDOM}};
  rob_uop_47_dst_value = _RAND_498[63:0];
  _RAND_499 = {2{`RANDOM}};
  rob_uop_47_src1_value = _RAND_499[63:0];
  _RAND_500 = {1{`RANDOM}};
  rob_uop_47_alu_sel = _RAND_500[4:0];
  _RAND_501 = {1{`RANDOM}};
  rob_uop_48_pc = _RAND_501[31:0];
  _RAND_502 = {1{`RANDOM}};
  rob_uop_48_inst = _RAND_502[31:0];
  _RAND_503 = {1{`RANDOM}};
  rob_uop_48_func_code = _RAND_503[6:0];
  _RAND_504 = {1{`RANDOM}};
  rob_uop_48_phy_dst = _RAND_504[6:0];
  _RAND_505 = {1{`RANDOM}};
  rob_uop_48_stale_dst = _RAND_505[6:0];
  _RAND_506 = {1{`RANDOM}};
  rob_uop_48_arch_dst = _RAND_506[4:0];
  _RAND_507 = {2{`RANDOM}};
  rob_uop_48_dst_value = _RAND_507[63:0];
  _RAND_508 = {2{`RANDOM}};
  rob_uop_48_src1_value = _RAND_508[63:0];
  _RAND_509 = {1{`RANDOM}};
  rob_uop_48_alu_sel = _RAND_509[4:0];
  _RAND_510 = {1{`RANDOM}};
  rob_uop_49_pc = _RAND_510[31:0];
  _RAND_511 = {1{`RANDOM}};
  rob_uop_49_inst = _RAND_511[31:0];
  _RAND_512 = {1{`RANDOM}};
  rob_uop_49_func_code = _RAND_512[6:0];
  _RAND_513 = {1{`RANDOM}};
  rob_uop_49_phy_dst = _RAND_513[6:0];
  _RAND_514 = {1{`RANDOM}};
  rob_uop_49_stale_dst = _RAND_514[6:0];
  _RAND_515 = {1{`RANDOM}};
  rob_uop_49_arch_dst = _RAND_515[4:0];
  _RAND_516 = {2{`RANDOM}};
  rob_uop_49_dst_value = _RAND_516[63:0];
  _RAND_517 = {2{`RANDOM}};
  rob_uop_49_src1_value = _RAND_517[63:0];
  _RAND_518 = {1{`RANDOM}};
  rob_uop_49_alu_sel = _RAND_518[4:0];
  _RAND_519 = {1{`RANDOM}};
  rob_uop_50_pc = _RAND_519[31:0];
  _RAND_520 = {1{`RANDOM}};
  rob_uop_50_inst = _RAND_520[31:0];
  _RAND_521 = {1{`RANDOM}};
  rob_uop_50_func_code = _RAND_521[6:0];
  _RAND_522 = {1{`RANDOM}};
  rob_uop_50_phy_dst = _RAND_522[6:0];
  _RAND_523 = {1{`RANDOM}};
  rob_uop_50_stale_dst = _RAND_523[6:0];
  _RAND_524 = {1{`RANDOM}};
  rob_uop_50_arch_dst = _RAND_524[4:0];
  _RAND_525 = {2{`RANDOM}};
  rob_uop_50_dst_value = _RAND_525[63:0];
  _RAND_526 = {2{`RANDOM}};
  rob_uop_50_src1_value = _RAND_526[63:0];
  _RAND_527 = {1{`RANDOM}};
  rob_uop_50_alu_sel = _RAND_527[4:0];
  _RAND_528 = {1{`RANDOM}};
  rob_uop_51_pc = _RAND_528[31:0];
  _RAND_529 = {1{`RANDOM}};
  rob_uop_51_inst = _RAND_529[31:0];
  _RAND_530 = {1{`RANDOM}};
  rob_uop_51_func_code = _RAND_530[6:0];
  _RAND_531 = {1{`RANDOM}};
  rob_uop_51_phy_dst = _RAND_531[6:0];
  _RAND_532 = {1{`RANDOM}};
  rob_uop_51_stale_dst = _RAND_532[6:0];
  _RAND_533 = {1{`RANDOM}};
  rob_uop_51_arch_dst = _RAND_533[4:0];
  _RAND_534 = {2{`RANDOM}};
  rob_uop_51_dst_value = _RAND_534[63:0];
  _RAND_535 = {2{`RANDOM}};
  rob_uop_51_src1_value = _RAND_535[63:0];
  _RAND_536 = {1{`RANDOM}};
  rob_uop_51_alu_sel = _RAND_536[4:0];
  _RAND_537 = {1{`RANDOM}};
  rob_uop_52_pc = _RAND_537[31:0];
  _RAND_538 = {1{`RANDOM}};
  rob_uop_52_inst = _RAND_538[31:0];
  _RAND_539 = {1{`RANDOM}};
  rob_uop_52_func_code = _RAND_539[6:0];
  _RAND_540 = {1{`RANDOM}};
  rob_uop_52_phy_dst = _RAND_540[6:0];
  _RAND_541 = {1{`RANDOM}};
  rob_uop_52_stale_dst = _RAND_541[6:0];
  _RAND_542 = {1{`RANDOM}};
  rob_uop_52_arch_dst = _RAND_542[4:0];
  _RAND_543 = {2{`RANDOM}};
  rob_uop_52_dst_value = _RAND_543[63:0];
  _RAND_544 = {2{`RANDOM}};
  rob_uop_52_src1_value = _RAND_544[63:0];
  _RAND_545 = {1{`RANDOM}};
  rob_uop_52_alu_sel = _RAND_545[4:0];
  _RAND_546 = {1{`RANDOM}};
  rob_uop_53_pc = _RAND_546[31:0];
  _RAND_547 = {1{`RANDOM}};
  rob_uop_53_inst = _RAND_547[31:0];
  _RAND_548 = {1{`RANDOM}};
  rob_uop_53_func_code = _RAND_548[6:0];
  _RAND_549 = {1{`RANDOM}};
  rob_uop_53_phy_dst = _RAND_549[6:0];
  _RAND_550 = {1{`RANDOM}};
  rob_uop_53_stale_dst = _RAND_550[6:0];
  _RAND_551 = {1{`RANDOM}};
  rob_uop_53_arch_dst = _RAND_551[4:0];
  _RAND_552 = {2{`RANDOM}};
  rob_uop_53_dst_value = _RAND_552[63:0];
  _RAND_553 = {2{`RANDOM}};
  rob_uop_53_src1_value = _RAND_553[63:0];
  _RAND_554 = {1{`RANDOM}};
  rob_uop_53_alu_sel = _RAND_554[4:0];
  _RAND_555 = {1{`RANDOM}};
  rob_uop_54_pc = _RAND_555[31:0];
  _RAND_556 = {1{`RANDOM}};
  rob_uop_54_inst = _RAND_556[31:0];
  _RAND_557 = {1{`RANDOM}};
  rob_uop_54_func_code = _RAND_557[6:0];
  _RAND_558 = {1{`RANDOM}};
  rob_uop_54_phy_dst = _RAND_558[6:0];
  _RAND_559 = {1{`RANDOM}};
  rob_uop_54_stale_dst = _RAND_559[6:0];
  _RAND_560 = {1{`RANDOM}};
  rob_uop_54_arch_dst = _RAND_560[4:0];
  _RAND_561 = {2{`RANDOM}};
  rob_uop_54_dst_value = _RAND_561[63:0];
  _RAND_562 = {2{`RANDOM}};
  rob_uop_54_src1_value = _RAND_562[63:0];
  _RAND_563 = {1{`RANDOM}};
  rob_uop_54_alu_sel = _RAND_563[4:0];
  _RAND_564 = {1{`RANDOM}};
  rob_uop_55_pc = _RAND_564[31:0];
  _RAND_565 = {1{`RANDOM}};
  rob_uop_55_inst = _RAND_565[31:0];
  _RAND_566 = {1{`RANDOM}};
  rob_uop_55_func_code = _RAND_566[6:0];
  _RAND_567 = {1{`RANDOM}};
  rob_uop_55_phy_dst = _RAND_567[6:0];
  _RAND_568 = {1{`RANDOM}};
  rob_uop_55_stale_dst = _RAND_568[6:0];
  _RAND_569 = {1{`RANDOM}};
  rob_uop_55_arch_dst = _RAND_569[4:0];
  _RAND_570 = {2{`RANDOM}};
  rob_uop_55_dst_value = _RAND_570[63:0];
  _RAND_571 = {2{`RANDOM}};
  rob_uop_55_src1_value = _RAND_571[63:0];
  _RAND_572 = {1{`RANDOM}};
  rob_uop_55_alu_sel = _RAND_572[4:0];
  _RAND_573 = {1{`RANDOM}};
  rob_uop_56_pc = _RAND_573[31:0];
  _RAND_574 = {1{`RANDOM}};
  rob_uop_56_inst = _RAND_574[31:0];
  _RAND_575 = {1{`RANDOM}};
  rob_uop_56_func_code = _RAND_575[6:0];
  _RAND_576 = {1{`RANDOM}};
  rob_uop_56_phy_dst = _RAND_576[6:0];
  _RAND_577 = {1{`RANDOM}};
  rob_uop_56_stale_dst = _RAND_577[6:0];
  _RAND_578 = {1{`RANDOM}};
  rob_uop_56_arch_dst = _RAND_578[4:0];
  _RAND_579 = {2{`RANDOM}};
  rob_uop_56_dst_value = _RAND_579[63:0];
  _RAND_580 = {2{`RANDOM}};
  rob_uop_56_src1_value = _RAND_580[63:0];
  _RAND_581 = {1{`RANDOM}};
  rob_uop_56_alu_sel = _RAND_581[4:0];
  _RAND_582 = {1{`RANDOM}};
  rob_uop_57_pc = _RAND_582[31:0];
  _RAND_583 = {1{`RANDOM}};
  rob_uop_57_inst = _RAND_583[31:0];
  _RAND_584 = {1{`RANDOM}};
  rob_uop_57_func_code = _RAND_584[6:0];
  _RAND_585 = {1{`RANDOM}};
  rob_uop_57_phy_dst = _RAND_585[6:0];
  _RAND_586 = {1{`RANDOM}};
  rob_uop_57_stale_dst = _RAND_586[6:0];
  _RAND_587 = {1{`RANDOM}};
  rob_uop_57_arch_dst = _RAND_587[4:0];
  _RAND_588 = {2{`RANDOM}};
  rob_uop_57_dst_value = _RAND_588[63:0];
  _RAND_589 = {2{`RANDOM}};
  rob_uop_57_src1_value = _RAND_589[63:0];
  _RAND_590 = {1{`RANDOM}};
  rob_uop_57_alu_sel = _RAND_590[4:0];
  _RAND_591 = {1{`RANDOM}};
  rob_uop_58_pc = _RAND_591[31:0];
  _RAND_592 = {1{`RANDOM}};
  rob_uop_58_inst = _RAND_592[31:0];
  _RAND_593 = {1{`RANDOM}};
  rob_uop_58_func_code = _RAND_593[6:0];
  _RAND_594 = {1{`RANDOM}};
  rob_uop_58_phy_dst = _RAND_594[6:0];
  _RAND_595 = {1{`RANDOM}};
  rob_uop_58_stale_dst = _RAND_595[6:0];
  _RAND_596 = {1{`RANDOM}};
  rob_uop_58_arch_dst = _RAND_596[4:0];
  _RAND_597 = {2{`RANDOM}};
  rob_uop_58_dst_value = _RAND_597[63:0];
  _RAND_598 = {2{`RANDOM}};
  rob_uop_58_src1_value = _RAND_598[63:0];
  _RAND_599 = {1{`RANDOM}};
  rob_uop_58_alu_sel = _RAND_599[4:0];
  _RAND_600 = {1{`RANDOM}};
  rob_uop_59_pc = _RAND_600[31:0];
  _RAND_601 = {1{`RANDOM}};
  rob_uop_59_inst = _RAND_601[31:0];
  _RAND_602 = {1{`RANDOM}};
  rob_uop_59_func_code = _RAND_602[6:0];
  _RAND_603 = {1{`RANDOM}};
  rob_uop_59_phy_dst = _RAND_603[6:0];
  _RAND_604 = {1{`RANDOM}};
  rob_uop_59_stale_dst = _RAND_604[6:0];
  _RAND_605 = {1{`RANDOM}};
  rob_uop_59_arch_dst = _RAND_605[4:0];
  _RAND_606 = {2{`RANDOM}};
  rob_uop_59_dst_value = _RAND_606[63:0];
  _RAND_607 = {2{`RANDOM}};
  rob_uop_59_src1_value = _RAND_607[63:0];
  _RAND_608 = {1{`RANDOM}};
  rob_uop_59_alu_sel = _RAND_608[4:0];
  _RAND_609 = {1{`RANDOM}};
  rob_uop_60_pc = _RAND_609[31:0];
  _RAND_610 = {1{`RANDOM}};
  rob_uop_60_inst = _RAND_610[31:0];
  _RAND_611 = {1{`RANDOM}};
  rob_uop_60_func_code = _RAND_611[6:0];
  _RAND_612 = {1{`RANDOM}};
  rob_uop_60_phy_dst = _RAND_612[6:0];
  _RAND_613 = {1{`RANDOM}};
  rob_uop_60_stale_dst = _RAND_613[6:0];
  _RAND_614 = {1{`RANDOM}};
  rob_uop_60_arch_dst = _RAND_614[4:0];
  _RAND_615 = {2{`RANDOM}};
  rob_uop_60_dst_value = _RAND_615[63:0];
  _RAND_616 = {2{`RANDOM}};
  rob_uop_60_src1_value = _RAND_616[63:0];
  _RAND_617 = {1{`RANDOM}};
  rob_uop_60_alu_sel = _RAND_617[4:0];
  _RAND_618 = {1{`RANDOM}};
  rob_uop_61_pc = _RAND_618[31:0];
  _RAND_619 = {1{`RANDOM}};
  rob_uop_61_inst = _RAND_619[31:0];
  _RAND_620 = {1{`RANDOM}};
  rob_uop_61_func_code = _RAND_620[6:0];
  _RAND_621 = {1{`RANDOM}};
  rob_uop_61_phy_dst = _RAND_621[6:0];
  _RAND_622 = {1{`RANDOM}};
  rob_uop_61_stale_dst = _RAND_622[6:0];
  _RAND_623 = {1{`RANDOM}};
  rob_uop_61_arch_dst = _RAND_623[4:0];
  _RAND_624 = {2{`RANDOM}};
  rob_uop_61_dst_value = _RAND_624[63:0];
  _RAND_625 = {2{`RANDOM}};
  rob_uop_61_src1_value = _RAND_625[63:0];
  _RAND_626 = {1{`RANDOM}};
  rob_uop_61_alu_sel = _RAND_626[4:0];
  _RAND_627 = {1{`RANDOM}};
  rob_uop_62_pc = _RAND_627[31:0];
  _RAND_628 = {1{`RANDOM}};
  rob_uop_62_inst = _RAND_628[31:0];
  _RAND_629 = {1{`RANDOM}};
  rob_uop_62_func_code = _RAND_629[6:0];
  _RAND_630 = {1{`RANDOM}};
  rob_uop_62_phy_dst = _RAND_630[6:0];
  _RAND_631 = {1{`RANDOM}};
  rob_uop_62_stale_dst = _RAND_631[6:0];
  _RAND_632 = {1{`RANDOM}};
  rob_uop_62_arch_dst = _RAND_632[4:0];
  _RAND_633 = {2{`RANDOM}};
  rob_uop_62_dst_value = _RAND_633[63:0];
  _RAND_634 = {2{`RANDOM}};
  rob_uop_62_src1_value = _RAND_634[63:0];
  _RAND_635 = {1{`RANDOM}};
  rob_uop_62_alu_sel = _RAND_635[4:0];
  _RAND_636 = {1{`RANDOM}};
  rob_uop_63_pc = _RAND_636[31:0];
  _RAND_637 = {1{`RANDOM}};
  rob_uop_63_inst = _RAND_637[31:0];
  _RAND_638 = {1{`RANDOM}};
  rob_uop_63_func_code = _RAND_638[6:0];
  _RAND_639 = {1{`RANDOM}};
  rob_uop_63_phy_dst = _RAND_639[6:0];
  _RAND_640 = {1{`RANDOM}};
  rob_uop_63_stale_dst = _RAND_640[6:0];
  _RAND_641 = {1{`RANDOM}};
  rob_uop_63_arch_dst = _RAND_641[4:0];
  _RAND_642 = {2{`RANDOM}};
  rob_uop_63_dst_value = _RAND_642[63:0];
  _RAND_643 = {2{`RANDOM}};
  rob_uop_63_src1_value = _RAND_643[63:0];
  _RAND_644 = {1{`RANDOM}};
  rob_uop_63_alu_sel = _RAND_644[4:0];
  _RAND_645 = {1{`RANDOM}};
  rob_done_0 = _RAND_645[0:0];
  _RAND_646 = {1{`RANDOM}};
  rob_done_1 = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  rob_done_2 = _RAND_647[0:0];
  _RAND_648 = {1{`RANDOM}};
  rob_done_3 = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  rob_done_4 = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  rob_done_5 = _RAND_650[0:0];
  _RAND_651 = {1{`RANDOM}};
  rob_done_6 = _RAND_651[0:0];
  _RAND_652 = {1{`RANDOM}};
  rob_done_7 = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  rob_done_8 = _RAND_653[0:0];
  _RAND_654 = {1{`RANDOM}};
  rob_done_9 = _RAND_654[0:0];
  _RAND_655 = {1{`RANDOM}};
  rob_done_10 = _RAND_655[0:0];
  _RAND_656 = {1{`RANDOM}};
  rob_done_11 = _RAND_656[0:0];
  _RAND_657 = {1{`RANDOM}};
  rob_done_12 = _RAND_657[0:0];
  _RAND_658 = {1{`RANDOM}};
  rob_done_13 = _RAND_658[0:0];
  _RAND_659 = {1{`RANDOM}};
  rob_done_14 = _RAND_659[0:0];
  _RAND_660 = {1{`RANDOM}};
  rob_done_15 = _RAND_660[0:0];
  _RAND_661 = {1{`RANDOM}};
  rob_done_16 = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  rob_done_17 = _RAND_662[0:0];
  _RAND_663 = {1{`RANDOM}};
  rob_done_18 = _RAND_663[0:0];
  _RAND_664 = {1{`RANDOM}};
  rob_done_19 = _RAND_664[0:0];
  _RAND_665 = {1{`RANDOM}};
  rob_done_20 = _RAND_665[0:0];
  _RAND_666 = {1{`RANDOM}};
  rob_done_21 = _RAND_666[0:0];
  _RAND_667 = {1{`RANDOM}};
  rob_done_22 = _RAND_667[0:0];
  _RAND_668 = {1{`RANDOM}};
  rob_done_23 = _RAND_668[0:0];
  _RAND_669 = {1{`RANDOM}};
  rob_done_24 = _RAND_669[0:0];
  _RAND_670 = {1{`RANDOM}};
  rob_done_25 = _RAND_670[0:0];
  _RAND_671 = {1{`RANDOM}};
  rob_done_26 = _RAND_671[0:0];
  _RAND_672 = {1{`RANDOM}};
  rob_done_27 = _RAND_672[0:0];
  _RAND_673 = {1{`RANDOM}};
  rob_done_28 = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  rob_done_29 = _RAND_674[0:0];
  _RAND_675 = {1{`RANDOM}};
  rob_done_30 = _RAND_675[0:0];
  _RAND_676 = {1{`RANDOM}};
  rob_done_31 = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  rob_done_32 = _RAND_677[0:0];
  _RAND_678 = {1{`RANDOM}};
  rob_done_33 = _RAND_678[0:0];
  _RAND_679 = {1{`RANDOM}};
  rob_done_34 = _RAND_679[0:0];
  _RAND_680 = {1{`RANDOM}};
  rob_done_35 = _RAND_680[0:0];
  _RAND_681 = {1{`RANDOM}};
  rob_done_36 = _RAND_681[0:0];
  _RAND_682 = {1{`RANDOM}};
  rob_done_37 = _RAND_682[0:0];
  _RAND_683 = {1{`RANDOM}};
  rob_done_38 = _RAND_683[0:0];
  _RAND_684 = {1{`RANDOM}};
  rob_done_39 = _RAND_684[0:0];
  _RAND_685 = {1{`RANDOM}};
  rob_done_40 = _RAND_685[0:0];
  _RAND_686 = {1{`RANDOM}};
  rob_done_41 = _RAND_686[0:0];
  _RAND_687 = {1{`RANDOM}};
  rob_done_42 = _RAND_687[0:0];
  _RAND_688 = {1{`RANDOM}};
  rob_done_43 = _RAND_688[0:0];
  _RAND_689 = {1{`RANDOM}};
  rob_done_44 = _RAND_689[0:0];
  _RAND_690 = {1{`RANDOM}};
  rob_done_45 = _RAND_690[0:0];
  _RAND_691 = {1{`RANDOM}};
  rob_done_46 = _RAND_691[0:0];
  _RAND_692 = {1{`RANDOM}};
  rob_done_47 = _RAND_692[0:0];
  _RAND_693 = {1{`RANDOM}};
  rob_done_48 = _RAND_693[0:0];
  _RAND_694 = {1{`RANDOM}};
  rob_done_49 = _RAND_694[0:0];
  _RAND_695 = {1{`RANDOM}};
  rob_done_50 = _RAND_695[0:0];
  _RAND_696 = {1{`RANDOM}};
  rob_done_51 = _RAND_696[0:0];
  _RAND_697 = {1{`RANDOM}};
  rob_done_52 = _RAND_697[0:0];
  _RAND_698 = {1{`RANDOM}};
  rob_done_53 = _RAND_698[0:0];
  _RAND_699 = {1{`RANDOM}};
  rob_done_54 = _RAND_699[0:0];
  _RAND_700 = {1{`RANDOM}};
  rob_done_55 = _RAND_700[0:0];
  _RAND_701 = {1{`RANDOM}};
  rob_done_56 = _RAND_701[0:0];
  _RAND_702 = {1{`RANDOM}};
  rob_done_57 = _RAND_702[0:0];
  _RAND_703 = {1{`RANDOM}};
  rob_done_58 = _RAND_703[0:0];
  _RAND_704 = {1{`RANDOM}};
  rob_done_59 = _RAND_704[0:0];
  _RAND_705 = {1{`RANDOM}};
  rob_done_60 = _RAND_705[0:0];
  _RAND_706 = {1{`RANDOM}};
  rob_done_61 = _RAND_706[0:0];
  _RAND_707 = {1{`RANDOM}};
  rob_done_62 = _RAND_707[0:0];
  _RAND_708 = {1{`RANDOM}};
  rob_done_63 = _RAND_708[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
